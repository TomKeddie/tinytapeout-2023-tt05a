module vga(
	       input  clk,
	       input  rst,
	       output r0,
	       output r1,
	       output r2,
	       output r3,
	       output g0,
	       output g1,
	       output g2,
	       output g3,
	       output b0,
	       output b1,
	       output b2,
	       output b3,
	       output hs,
	       output vs
	       );

  localparam	  h_visible    = 640;
  localparam	  h_frontporch = 640 + 16;
  localparam	  h_sync       = 640 + 16 + 96;
  localparam	  h_backporch  = 640 + 16 + 96 + 47;

  // while h_sync is being sent, vertical counts h_sync pulses, for
  // porch and sync, it counts clocks
  localparam	  v_visible    = 480;
  localparam	  v_frontporch = 480 + 22;
  localparam	  v_sync       = 480 + 22 + 3;
  localparam	  v_backporch = 480 + 22 + 3 + 1;

  localparam smile001  = 59'b00000000000000000000000000000000000000000000000000010000000;
  localparam smile002  = 59'b00000000000000000000000000000000000000000000000000111000000;
  localparam smile003  = 59'b00000000000000000000000000000000000000000000000000111110000;
  localparam smile004  = 59'b00000000000000000000000000000000000000000000000001111111000;
  localparam smile005  = 59'b00000000000000000000000000000000000000000000000011111111100;
  localparam smile006  = 59'b00000000000000000000000000000000000000000000000111111111110;
  localparam smile007  = 59'b00000000000000000000000000000000000000000000000111111111110;
  localparam smile008  = 59'b00000000000000000000000000000000000000000000001111111111100;
  localparam smile009  = 59'b00000000000000000000000000000000000000000000011111111111100;
  localparam smile010  = 59'b00000000000000000000000000000000000000000000011111111111000;
  localparam smile011  = 59'b00000000000000000000000000000000000000000000111111111110000;
  localparam smile012  = 59'b00000000000000000000000000000000000000000001111111111110000;
  localparam smile013  = 59'b00000000000000000000000000000000000000000001111111111100000;
  localparam smile014  = 59'b00000000000000000000000000000000000000000011111111111100000;
  localparam smile015  = 59'b00000000000000000000000000000000000000000011111111111000000;
  localparam smile016  = 59'b00000000000000000000000000000000000000000111111111110000000;
  localparam smile017  = 59'b00000000000000000000000000000000000000000111111111110000000;
  localparam smile018  = 59'b00000000000000000000000000000000000000001111111111100000000;
  localparam smile019  = 59'b00000000000000000000000000000000000000001111111111100000000;
  localparam smile020  = 59'b00000000000000000000000000000000000000011111111111000000000;
  localparam smile021  = 59'b00000000000000000000000000000000000000011111111111000000000;
  localparam smile022  = 59'b00000000000000000000000000000000000000111111111111000000000;
  localparam smile023  = 59'b00000000000000000000000000000000000000111111111110000000000;
  localparam smile024  = 59'b00000000000000000000000000000000000001111111111110000000000;
  localparam smile025  = 59'b00000000000000000000000000000000000001111111111100000000000;
  localparam smile026  = 59'b00000000000000000000000000000000000001111111111100000000000;
  localparam smile027  = 59'b00000000000000000000000000000000000011111111111100000000000;
  localparam smile028  = 59'b00000111111100000000000000000000000011111111111000000000000;
  localparam smile029  = 59'b00011111111111000000000000000000000011111111111000000000000;
  localparam smile030  = 59'b00111111111111100000000000000000000111111111111000000000000;
  localparam smile031  = 59'b01111111111111110000000000000000000111111111110000000000000;
  localparam smile032  = 59'b11111111111111111000000000000000000111111111110000000000000;
  localparam smile033  = 59'b11111111111111111000000000000000000111111111110000000000000;
  localparam smile034  = 59'b11111111111111111000000000000000001111111111110000000000000;
  localparam smile035  = 59'b11111111111111111100000000000000001111111111100000000000000;
  localparam smile036  = 59'b11111111111111111100000000000000001111111111100000000000000;
  localparam smile037  = 59'b11111111111111111100000000000000001111111111100000000000000;
  localparam smile038  = 59'b11111111111111111000000000000000001111111111100000000000000;
  localparam smile039  = 59'b11111111111111111000000000000000001111111111100000000000000;
  localparam smile040  = 59'b01111111111111111000000000000000011111111111000000000000000;
  localparam smile041  = 59'b01111111111111110000000000000000011111111111000000000000000;
  localparam smile042  = 59'b00111111111111100000000000000000011111111111000000000000000;
  localparam smile043  = 59'b00011111111111000000000000000000011111111111000000000000000;
  localparam smile044  = 59'b00000111111100000000000000000000011111111111000000000000000;
  localparam smile045  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile046  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile047  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile048  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile049  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile050  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile051  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile052  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile053  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile054  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile055  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile056  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile057  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile058  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile059  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile060  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile061  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile062  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile063  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile064  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile065  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile066  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile067  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile068  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile069  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile070  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile071  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile072  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile073  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile074  = 59'b00000000000000000000000000000000011111111111100000000000000;
  localparam smile075  = 59'b00000000000000000000000000000000001111111111100000000000000;
  localparam smile076  = 59'b00000000000000000000000000000000001111111111100000000000000;
  localparam smile077  = 59'b00000001110000000000000000000000001111111111100000000000000;
  localparam smile078  = 59'b00001111111110000000000000000000001111111111100000000000000;
  localparam smile079  = 59'b00011111111111100000000000000000001111111111110000000000000;
  localparam smile080  = 59'b00111111111111110000000000000000000111111111110000000000000;
  localparam smile081  = 59'b01111111111111110000000000000000000111111111110000000000000;
  localparam smile082  = 59'b11111111111111111000000000000000000111111111111000000000000;
  localparam smile083  = 59'b11111111111111111000000000000000000111111111111000000000000;
  localparam smile084  = 59'b11111111111111111000000000000000000011111111111000000000000;
  localparam smile085  = 59'b11111111111111111100000000000000000011111111111100000000000;
  localparam smile086  = 59'b11111111111111111100000000000000000011111111111100000000000;
  localparam smile087  = 59'b11111111111111111000000000000000000001111111111100000000000;
  localparam smile088  = 59'b11111111111111111000000000000000000001111111111110000000000;
  localparam smile089  = 59'b11111111111111111000000000000000000001111111111110000000000;
  localparam smile090  = 59'b01111111111111110000000000000000000000111111111110000000000;
  localparam smile091  = 59'b00111111111111110000000000000000000000111111111111000000000;
  localparam smile092  = 59'b00111111111111100000000000000000000000111111111111000000000;
  localparam smile093  = 59'b00001111111110000000000000000000000000011111111111100000000;
  localparam smile094  = 59'b00000011111000000000000000000000000000011111111111100000000;
  localparam smile095  = 59'b00000000000000000000000000000000000000001111111111110000000;
  localparam smile096  = 59'b00000000000000000000000000000000000000001111111111110000000;
  localparam smile097  = 59'b00000000000000000000000000000000000000000111111111111000000;
  localparam smile098  = 59'b00000000000000000000000000000000000000000111111111111000000;
  localparam smile099  = 59'b00000000000000000000000000000000000000000011111111111100000;
  localparam smile100  = 59'b00000000000000000000000000000000000000000001111111111110000;
  localparam smile101  = 59'b00000000000000000000000000000000000000000001111111111110000;
  localparam smile102  = 59'b00000000000000000000000000000000000000000000111111111111000;
  localparam smile103  = 59'b00000000000000000000000000000000000000000000111111111111000;
  localparam smile104  = 59'b00000000000000000000000000000000000000000000011111111111100;
  localparam smile105  = 59'b00000000000000000000000000000000000000000000001111111111110;
  localparam smile106  = 59'b00000000000000000000000000000000000000000000000111111111110;
  localparam smile107  = 59'b00000000000000000000000000000000000000000000000111111111111;
  localparam smile108  = 59'b00000000000000000000000000000000000000000000000011111111110;
  localparam smile109  = 59'b00000000000000000000000000000000000000000000000001111111100;
  localparam smile110  = 59'b00000000000000000000000000000000000000000000000000111111000;
  localparam smile111  = 59'b00000000000000000000000000000000000000000000000000011110000;
  localparam smile112  = 59'b00000000000000000000000000000000000000000000000000011000000;


  localparam words01  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000;
  localparam words02  = 506'b11110000000000011100000000000000000000000000000000000000000000000000000000000000011110000000000000001111111110000000111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000;
  localparam words03  = 506'b01110000000000111100000000000000000000000000000000000000000000000000000000000000011111000000000000111111111111000000111000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words04  = 506'b01111000000001111000000000000000000000000000000000000000000000000000000000000000111111000000000001111111111111000000111000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000;
  localparam words05  = 506'b00111100000001110000000000000000000000000000000000000000000000000000000000000000111111100000000011111100001111000000111000000011111100000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000;
  localparam words06  = 506'b00011100000011110000000000000000000000000000000000000000000000000000000000000000111011100000000011110000000000000000111000000111110000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000;
  localparam words07  = 506'b00011110000111100000000000000000000000000000000000000000000000000000000000000001111011100000000011100000000000000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000;
  localparam words08  = 506'b00001111000111000000111111100000001111000000011110000111100111110000000000000001110011110000000011100000000000000000111000001111000000000000000000000000000111100111110001111111100000000111100111111000000000000000000111000011110011111100000011111111110000000111111100000000000000000001111111100000000000000000011110011111100000001111001111100000111111100000001111001111110000000011100000000111111100000001111001111100000111111000000000000000000111000111111111100000000000000000000000000000000000000000000000;
  localparam words09  = 506'b00000111001111000011111111110000001111000000011110000111111111110000000000000011110001110000000011110000000000000000111000001111000000000000000000000000000111111111110011111111111000000111111111111100000000000000000111000011111111111110000011111111110000011111111110000000000000000011111111111000000000000000011111111111110000001111111111100011111111110000001111111111111000000011100000011111111111000001111111111111001111111100000000000000000111000111111111100000000000000000000000000000000000000000000000;
  localparam words10  = 506'b00000111111110000111111111111000001111000000011110000111111111110000000000000011110001110000000011111000000000000000111000001110000000000000000000000000000111111111110011111111111100000111111111111110000000000000000111000011111111111111000011111111110000111111111111000000000000000011111111111100000000000000011111111111111000001111111111100111111111111000001111111111111100000011100000111111111111100001111111111111011111111110000000000000000111000111111111100000000000000000000000000000000000000000000000;
  localparam words11  = 506'b00000011111100001111110001111100001111000000011110000111111100000000000000000011100001111000000001111111100000000000111000001110000000000000000000000000000111111100000011100001111100000111111100111110000000000000000111000011111110011111000001111000000001111110001111100000000000000011100001111100000000000000011111110011111100001111111000001111110001111100001111111001111110000011100000111110001111100001111110001111111100011110000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words12  = 506'b00000001111100001111000000111100001111000000011110000111110000000000000000000111100000111000000000111111111100000000111000011110000000000000000000000000000111110000000000000000011110000111110000001111000000000000000111000011111000000111100001111000000001111000000111100000000000000000000000011110000000000000011111000000111100001111100000001111000000111100001111100000011110000011100001111000000011110001111100000011110000001111000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words13  = 506'b00000001111000001110000000011110001111000000011110000111100000000000000000000111000000111100000000011111111111000000111000011110000000000000000000000000000111100000000000000000001110000111100000001111000000000000000111000011110000000111100001111000000001110000000011110000000000000000000000001110000000000000011110000000011100001111000000001110000000011110001111000000001110000011100001110000000001110001111000000011110000000111000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words14  = 506'b00000001111000011110000000011110001111000000011110000111100000000000000000000111000000111100000000000001111111100000111000001110000000000000000000000000000111100000000000111111111110000111100000001111000000000000000111000011110000000111100001111000000011110000000011110000000000000000111111111110000000000000011110000000011110001111000000011110000000011110001111000000001111000011100001111111111111110001111000000011100000000111000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words15  = 506'b00000001111000011110000000001110001111000000011110000111100000000000000000001111000000011100000000000000000111100000111000001110000000000000000000000000000111100000000011111111111110000111100000001111000000000000000111000011110000000111100001111000000011110000000001110000000000000011111111111110000000000000011110000000011110001111000000011110000000001110001111000000001111000011100011111111111111110001111000000011100000000111000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words16  = 506'b00000001111000011110000000001110001111000000011110000111100000000000000000001111111111111110000000000000000011110000111000001111000000000000000000000000000111100000000111111111111110000111100000001111000000000000000111000011110000000111100001111000000011110000000001110000000000000111111111111110000000000000011110000000011110001111000000011110000000001110001111000000001111000011100011111111111111110001111000000011100000000111000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words17  = 506'b00000001111000011110000000011110001111000000011110000111100000000000000000011111111111111110000000000000000011110000111000001111000000000000000000000000000111100000000111110000001110000111100000001111000000000000000111000011110000000111100001111000000011110000000011110000000000000111110000001110000000000000011110000000011110001111000000011110000000011110001111000000001111000011100011110000000000000001111000000011100000000111000000000000000111000011110000000000000000000000000000000000000000000000000000;
  localparam words18  = 506'b00000001111000001110000000011110001111000000011110000111100000000000000000011111111111111110000000000000000011110000111000000111100000000000000000000000000111100000000111000000011110000111100000001111000000000000000111000011110000000111100000111000000001110000000011110000000000000111000000011110000000000000011110000000011100001111000000001110000000011110001111000000001110000011100001110000000000000001111000000011100000000111000000000000000111000001110000000000000000000000000000000000000000000000000000;
  localparam words19  = 506'b00000001111000001111000000111100001111000000111110000111100000000000000000011100000000001111000000000000000111100000111000000111110000000000110000000000000111100000000111000000011110000111100000001111000000000000000111000011110000000111100000111000000001111000000111100000000000000111000000011110000000000000011111000000111100001111000000001111000000111100001111100000011110000011100001111000000000110001111000000011100000000111000000000000000111000001110000000000000000000000000000000000000000000000000000;
  localparam words20  = 506'b00000001111000001111110001111100000111110001111110000111100000000000000000111100000000000111000011110000011111100000111000000011111100000111110000000000000111100000000111100001111110000111100000001111000000000000000111000011110000000111100000111100000001111110001111100000000000000111100001111110000000000000011111110001111100001111000000001111110001111100001111111000111110000011100000111110000111110001111000000011100000000111000000000000000111000001111000000000000000000000000000000000000000000000000000;
  localparam words21  = 506'b00000001111000000111111111111000000111111111111110000111100000000000000000111100000000000111100011111111111111000000111000000001111111111111110000000000000111100000000111111111111110000111100000001111000000000000000111000011110000000111100000111111110000111111111111000000000000000111111111111110000000000000011111111111111000001111000000000111111111111000001111111111111100000011100000111111111111110001111000000011100000000111000000000000000111000001111111100000000000000000000000000000000000000000000000;
  localparam words22  = 506'b00000001111000000011111111110000000011111111111110000111100000000000000000111000000000000111100011111111111111000000111000000000111111111111100000000000000111100000000011111111101110000111100000001111000000000000000111000011110000000111100000111111110000011111111110000000000000000011111111101110000000000000011111111111110000001111000000000011111111110000001111111111111000000011100000011111111111100001111000000011100000000111000000000000000111000001111111100000000000000000000000000000000000000000000000;
  localparam words23  = 506'b00000001111000000000111111100000000001111110011110000111100000000000000001111000000000000011100001111111111100000000111000000000001111111110000000000000000111100000000001111111001110000111100000001111000000000000000111000011110000000111100000001111110000000111111100000000000000000001111111001110000000000000011110011111100000001111000000000000111111100000001111001111110000000011100000000111111110000001111000000011100000000111000000000000000111000000011111100000000000000000000000000000000000000000000000;
  localparam words24  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words25  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words26  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words27  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words28  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words29  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words30  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words31  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000011100000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words32  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000011100001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words33  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000011100001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words34  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000011100001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words35  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000011100001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words36  = 506'b00000000000000000000000000000000000000000000000000000000111000000000000000111100000000000000000000000011100001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
  localparam words37  = 506'b00000011111111000000001111111000000011110000000111100000111000000011111100111100001111001111110000000011100011111111110000000000000111100111111000000000111111110000000011110011111100000000001111110011110000011100000000111111100000000000000000000000000000111111110000000011110011111100000000001111110011110000000000000011110011111100000000000111111100000011100000011110000001110000000000000001110001111111111000000000000011110011111100000000000111111100000000000111111100000000001111110011110000001111111110;
  localparam words38  = 506'b00001111111111100000111111111100000011110000000111100000111000000111111111111100001111111111111000000011100011111111110000000000000111111111111100000001111111111100000011111111111110000000011111111111110000011100000011111111111000000000000000000000000001111111111100000011111111111110000000011111111111110000000000000011111111111110000000011111111110000011110000011111000001110000000000000001110001111111111000000000000011111111111110000000011111111111000000011111111111000000011111111111110000011111111111;
  localparam words39  = 506'b00011111111111100001111111111110000011110000000111100000111000001111111111111100001111111111111100000000000011111111110000000000000111111111111110000001111111111110000011111111111111000000111111111111110000011100000111111111111100000000000000000000000001111111111110000011111111111111000000111111111111110000000000000011111111111111000000111111111111000001110000011111000001110000000000000001110001111111111000000000000011111111111111000000111111111111100000111111111111100000111111111111110000111111111111;
  localparam words40  = 506'b00011111000011100011111100011111000011110000000111100000111000011111100011111100001111111001111100000000000001111000000000000000000111111100111110000001110000111110000011111110011111000001111110001111110000011100000111110001111100000000000000000000000001110000111110000011111110011111000001111110001111110000000000000011111110011111000001111110001111100001110000111111000011110000000000000001110000111100000000000000000011111110011111000000111110001111100000111110001111100001111110001111110000111100000111;
  localparam words41  = 506'b00111100000000000011110000001111000011110000000111100000111000011110000001111100001111100000011110000000000001111000000000000000000111110000001111000000000000001111000011111000000111100001111000000111110000011100001111000000011110000000000000000000000000000000001111000011111000000111100001111000000111110000000000000011111000000111100001111000000111100001110000111111000011100000000000000001110000111100000000000000000011111000000111100001111000000011110001111000000011110001111000000111110001111000000000;
  localparam words42  = 506'b00111000000000000011100000000111100011110000000111100000111000011100000000111100001111000000011110000000000001111000000000000000000111100000001111000000000000000111000011110000000111100001110000000011110000011100001110000000001110000000000000000000000000000000000111000011110000000111100001110000000011110000000000000011110000000111100001110000000011110001111000111011100011100000000000000001110000111100000000000000000011110000000111100001110000000001110001110000000001110001110000000011110000111000000000;
  localparam words43  = 506'b01111000000000000111100000000111100011110000000111100000111000111100000000111100001111000000011110000000000001111000000000000000000111100000001111000000011111111111000011110000000111100011110000000011110000011100001111111111111110000000000000000000000000011111111111000011110000000111100011110000000011110000000000000011110000000111100011110000000011110000111000111011100011100000000000000001110000111100000000000000000011110000000111100001111111111111110001111111111111110011110000000011110000111111100000;
  localparam words44  = 506'b01111000000000000111100000000011100011110000000111100000111000111100000000111100001111000000011110000000000001111000000000000000000111100000001111000001111111111111000011110000000111100011110000000011110000011100011111111111111110000000000000000000000001111111111111000011110000000111100011110000000011110000000000000011110000000111100011110000000001110000111001110011100111100000000000000001110000111100000000000000000011110000000111100011111111111111110011111111111111110011110000000011110000011111111100;
  localparam words45  = 506'b01111000000000000111100000000011100011110000000111100000111000111100000000111100001111000000011110000000000001111000000000000000000111100000001111000011111111111111000011110000000111100011110000000011110000011100011111111111111110000000000000000000000011111111111111000011110000000111100011110000000011110000000000000011110000000111100011110000000001110000111101110001100111000000000000000001110000111100000000000000000011110000000111100011111111111111110011111111111111110011110000000011110000000011111110;
  localparam words46  = 506'b01111000000000000111100000000111100011110000000111100000111000111100000000111100001111000000011110000000000001111000000000000000000111100000001111000011111000000111000011110000000111100011110000000011110000011100011110000000000000000000000000000000000011111000000111000011110000000111100011110000000011110000000000000011110000000111100011110000000011110000011101110001110111000000000000000001110000111100000000000000000011110000000111100011110000000000000011110000000000000011110000000011110000000000001111;
  localparam words47  = 506'b00111000000000000011100000000111100011110000000111100000111000011100000000111100001111000000011110000000000000111000000000000000000111100000001111000011100000001111000011110000000111100001110000000011110000011100001110000000000000000000000000000000000011100000001111000011110000000111100001110000000011110000000000000011110000000111100001110000000011110000011101110001111111000000000000000001110000011100000000000000000011110000000111100001110000000000000001110000000000000001110000000011110000000000000111;
  localparam words48  = 506'b00111100000000000011110000001111000011110000001111100000111000011110000001111100001111000000011110000000000000111000000000000000000111100000001111000011100000001111000011110000000111100001111000000111110000011100001111000000000110000000000000000000000011100000001111000011110000000111100001111000000111110000000000000011110000000111100001111000000111100000011111100001111110000000000000000001110000011100000000000000000011110000000111100001111000000000110001111000000000110001111000000111110001100000000111;
  localparam words49  = 506'b00011111000011100011111100011111000001111100011111100000111000011111100011111100001111000000011110000000000000111100000000000000000111100000001111000011110000111111000011110000000111100001111110001111110000011100000111110000111110000111100000000000000011110000111111000011110000000111100001111110001111110000000000000011110000000111100001111110001111100000011111100000111110000000000000000001110000011110000000000000000011110000000111100000111110000111110000111110000111110001111110001111110001111100011111;
  localparam words50  = 506'b00011111111111100001111111111110000001111111111111100000111000001111111111111100001111000000011110000000000000111111110000000000000111100000001111000011111111111111000011110000000111100000111111111111110000011100000111111111111110000111100000000000000011111111111111000011110000000111100000111111111111110000000000000011110000000111100000111111111111000000001111100000111110000000000000000001110000011111111000000000000011110000000111100000111111111111110000111111111111110000111111111111110001111111111111;
  localparam words51  = 506'b00001111111111100000111111111100000000111111111111100000111000000111111111111100001111000000011110000000000000111111110000000000000111100000001111000001111111110111000011110000000111100000011111111111110000011100000011111111111100000111100000000000000001111111110111000011110000000111100000011111111111110000000000000011110000000111100000011111111110000000001111000000111110000000000000000001110000011111111000000000000011110000000111100000011111111111100000011111111111100000011111111111110000111111111110;
  localparam words52  = 506'b00000011111111000000001111111000000000011111100111100000111000000011111110111100001111000000011110000000000000001111110000000000000111100000001111000000111111100111000011110000000111100000001111111011110000011100000000111111110000000111000000000000000000111111100111000011110000000111100000001111111011110000000000000011110000000111100000000111111100000000001111000000111100000000000000000001110000000111111000000000000011110000000111100000000111111110000000000111111110000000001111111011110000001111111000;
  localparam words53  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words54  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words55  = 506'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words56  = 506'b00111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words57  = 506'b00111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words58  = 506'b00111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words59  = 506'b00111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words60  = 506'b00111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words61  = 506'b01111111111000000011111110000000000000000011110011111000001111111000000000111111111000011111111110000011111111000000001111001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words62  = 506'b01111111111000001111111111000000000000000011111111111000111111111110000001111111111100011111111110000111111111110000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words63  = 506'b01111111111000011111111111100000000000000011111111111001111111111111000011111111111100011111111110000111111111111000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words64  = 506'b00111100000000111111000111110000000000000011111110000001111100011111000011110000011100001111000000000111000011111000001111111000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words65  = 506'b00111100000000111100000011110000000000000011111000000011110000000111100111100000000000001111000000000000000000111100001111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words66  = 506'b00111100000000111000000001111000000000000011110000000011100000000011100011100000000000001111000000000000000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words67  = 506'b00111100000001111000000001111000000000000011110000000011111111111111100011111110000000001111000000000001111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words68  = 506'b00111100000001111000000000111000000000000011110000000111111111111111100001111111110000001111000000000111111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words69  = 506'b00111100000001111000000000111000000000000011110000000111111111111111100000001111111000001111000000001111111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words70  = 506'b00111100000001111000000001111000000000000011110000000111100000000000000000000000111100001111000000001111100000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words71  = 506'b00011100000000111000000001111000000000000011110000000011100000000000000000000000011100000111000000001110000000111100001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words72  = 506'b00011100000000111100000011110000000000000011110000000011110000000001100110000000011100000111000000001110000000111100001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words73  = 506'b00011110000000111111000111110000000000000011110000000001111100001111100111110001111100000111100000001111000011111100001111000000000111100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words74  = 506'b00011111111000011111111111100000000000000011110000000001111111111111100111111111111100000111111110001111111111111100001111000000000111111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words75  = 506'b00011111111000001111111111000000000000000011110000000000111111111111000011111111111000000111111110000111111111011100001111000000000111111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words76  = 506'b00000111111000000011111110000000000000000011110000000000001111111100000000111111100000000001111110000011111110011100001111000000000001111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  

  wire            blank;
  reg             blank_h;
  reg             blank_v;

  assign blank = (blank_h | blank_v);

  // 2^10  = 1024
  reg [9:0]       count_h;
  // 2^15 = 32768
  reg [14:0]      count_v;

  wire            red;
  wire            grn;
  reg             blu;
  reg             wht;
  reg             hs_out;
  reg             vs_out;

  reg [3:0]       fb[3:0];

  assign r0 = red;
  assign r1 = red;
  assign r2 = red;
  assign r3 = red;
  assign b0 = blu;
  assign b1 = blu;
  assign b2 = blu;
  assign b3 = blu;
  assign g0 = grn;
  assign g1 = grn;
  assign g2 = grn;
  assign g3 = grn;
  assign hs = !hs_out;
  assign vs = !vs_out;

  assign red = wht;
  assign grn = wht;

  always @ (blank) begin
    if (blank) begin
      blu <= 1'b0;
      wht <= 1'b0;
    end else begin
      blu <= 1'b1;
      if (count_v > 99 && count_v < 211 && count_h > 80 && count_h < 140) begin
        case(count_v-99)
          1 : wht <= smile001[140-count_h];
          2 : wht <= smile002[140-count_h];
          3 : wht <= smile003[140-count_h];
          4 : wht <= smile004[140-count_h];
          5 : wht <= smile005[140-count_h];
          6 : wht <= smile006[140-count_h];
          7 : wht <= smile007[140-count_h];
          8 : wht <= smile008[140-count_h];
          9 : wht <= smile009[140-count_h];
          10 : wht <= smile010[140-count_h];
          11 : wht <= smile011[140-count_h];
          12 : wht <= smile012[140-count_h];
          13 : wht <= smile013[140-count_h];
          14 : wht <= smile014[140-count_h];
          15 : wht <= smile015[140-count_h];
          16 : wht <= smile016[140-count_h];
          17 : wht <= smile017[140-count_h];
          18 : wht <= smile018[140-count_h];
          19 : wht <= smile019[140-count_h];
          20 : wht <= smile020[140-count_h];
          21 : wht <= smile021[140-count_h];
          22 : wht <= smile022[140-count_h];
          23 : wht <= smile023[140-count_h];
          24 : wht <= smile024[140-count_h];
          25 : wht <= smile025[140-count_h];
          26 : wht <= smile026[140-count_h];
          27 : wht <= smile027[140-count_h];
          28 : wht <= smile028[140-count_h];
          80 : wht <= smile029[140-count_h];
          30 : wht <= smile030[140-count_h];
          31 : wht <= smile031[140-count_h];
          32 : wht <= smile032[140-count_h];
          33 : wht <= smile033[140-count_h];
          34 : wht <= smile034[140-count_h];
          35 : wht <= smile035[140-count_h];
          36 : wht <= smile036[140-count_h];
          37 : wht <= smile037[140-count_h];
          38 : wht <= smile038[140-count_h];
          39 : wht <= smile039[140-count_h];
          40 : wht <= smile040[140-count_h];
          41 : wht <= smile041[140-count_h];
          42 : wht <= smile042[140-count_h];
          43 : wht <= smile043[140-count_h];
          44 : wht <= smile044[140-count_h];
          45 : wht <= smile045[140-count_h];
          46 : wht <= smile046[140-count_h];
          47 : wht <= smile047[140-count_h];
          48 : wht <= smile048[140-count_h];
          49 : wht <= smile049[140-count_h];
          50 : wht <= smile050[140-count_h];
          51 : wht <= smile051[140-count_h];
          52 : wht <= smile052[140-count_h];
          53 : wht <= smile053[140-count_h];
          54 : wht <= smile054[140-count_h];
          55 : wht <= smile055[140-count_h];
          56 : wht <= smile056[140-count_h];
          57 : wht <= smile057[140-count_h];
          58 : wht <= smile058[140-count_h];
          59 : wht <= smile059[140-count_h];
          60 : wht <= smile060[140-count_h];
          61 : wht <= smile061[140-count_h];
          62 : wht <= smile062[140-count_h];
          63 : wht <= smile063[140-count_h];
          64 : wht <= smile064[140-count_h];
          65 : wht <= smile065[140-count_h];
          66 : wht <= smile066[140-count_h];
          67 : wht <= smile067[140-count_h];
          68 : wht <= smile068[140-count_h];
          69 : wht <= smile069[140-count_h];
          70 : wht <= smile070[140-count_h];
          71 : wht <= smile071[140-count_h];
          72 : wht <= smile072[140-count_h];
          73 : wht <= smile073[140-count_h];
          74 : wht <= smile074[140-count_h];
          75 : wht <= smile075[140-count_h];
          76 : wht <= smile076[140-count_h];
          77 : wht <= smile077[140-count_h];
          78 : wht <= smile078[140-count_h];
          79 : wht <= smile079[140-count_h];
          80 : wht <= smile080[140-count_h];
          81 : wht <= smile081[140-count_h];
          82 : wht <= smile082[140-count_h];
          83 : wht <= smile083[140-count_h];
          84 : wht <= smile084[140-count_h];
          85 : wht <= smile085[140-count_h];
          86 : wht <= smile086[140-count_h];
          87 : wht <= smile087[140-count_h];
          88 : wht <= smile088[140-count_h];
          89 : wht <= smile089[140-count_h];
          90 : wht <= smile090[140-count_h];
          91 : wht <= smile091[140-count_h];
          92 : wht <= smile092[140-count_h];
          93 : wht <= smile093[140-count_h];
          94 : wht <= smile094[140-count_h];
          95 : wht <= smile095[140-count_h];
          96 : wht <= smile096[140-count_h];
          97 : wht <= smile097[140-count_h];
          98 : wht <= smile098[140-count_h];
          99 : wht <= smile099[140-count_h];
          100 : wht <= smile100[140-count_h];
          101 : wht <= smile101[140-count_h];
          102 : wht <= smile102[140-count_h];
          103 : wht <= smile103[140-count_h];
          104 : wht <= smile104[140-count_h];
          105 : wht <= smile105[140-count_h];
          106 : wht <= smile106[140-count_h];
          107 : wht <= smile107[140-count_h];
          108 : wht <= smile108[140-count_h];
          109 : wht <= smile109[140-count_h];
          110 : wht <= smile110[140-count_h];
          111 : wht <= smile111[140-count_h];
          112 : wht <= smile112[140-count_h];
          default: wht <= 1'b0;
        endcase
      end else if (count_v > 299 && count_v < 376 && count_h > 40 && count_h < 546) begin
        case(count_v-299)
          1 : wht  <= words01[546-count_h];
          2 : wht  <= words02[546-count_h];
          3 : wht  <= words03[546-count_h];
          4 : wht  <= words04[546-count_h];
          5 : wht  <= words05[546-count_h];
          6 : wht  <= words06[546-count_h];
          7 : wht  <= words07[546-count_h];
          8 : wht  <= words08[546-count_h];
          9 : wht  <= words09[546-count_h];
          10 : wht <= words10[546-count_h];
          11 : wht <= words11[546-count_h];
          12 : wht <= words12[546-count_h];
          13 : wht <= words13[546-count_h];
          14 : wht <= words14[546-count_h];
          15 : wht <= words15[546-count_h];
          16 : wht <= words16[546-count_h];
          17 : wht <= words17[546-count_h];
          18 : wht <= words18[546-count_h];
          19 : wht <= words19[546-count_h];
          20 : wht <= words20[546-count_h];
          21 : wht <= words21[546-count_h];
          22 : wht <= words22[546-count_h];
          23 : wht <= words23[546-count_h];
          24 : wht <= words24[546-count_h];
          25 : wht <= words25[546-count_h];
          26 : wht <= words26[546-count_h];
          27 : wht <= words27[546-count_h];
          28 : wht <= words28[546-count_h];
          29 : wht <= words29[546-count_h];
          30 : wht <= words30[546-count_h];
          31 : wht <= words31[546-count_h];
          32 : wht <= words32[546-count_h];
          33 : wht <= words33[546-count_h];
          34 : wht <= words34[546-count_h];
          35 : wht <= words35[546-count_h];
          36 : wht <= words36[546-count_h];
          37 : wht <= words37[546-count_h];
          38 : wht <= words38[546-count_h];
          39 : wht <= words39[546-count_h];
          40 : wht <= words40[546-count_h];
          41 : wht <= words41[546-count_h];
          42 : wht <= words42[546-count_h];
          43 : wht <= words43[546-count_h];
          44 : wht <= words44[546-count_h];
          45 : wht <= words45[546-count_h];
          46 : wht <= words46[546-count_h];
          47 : wht <= words47[546-count_h];
          48 : wht <= words48[546-count_h];
          49 : wht <= words49[546-count_h];
          50 : wht <= words50[546-count_h];
          51 : wht <= words51[546-count_h];
          52 : wht <= words52[546-count_h];
          53 : wht <= words53[546-count_h];
          54 : wht <= words54[546-count_h];
          55 : wht <= words55[546-count_h];
          56 : wht <= words56[546-count_h];
          57 : wht <= words57[546-count_h];
          58 : wht <= words58[546-count_h];
          59 : wht <= words59[546-count_h];
          60 : wht <= words60[546-count_h];
          61 : wht <= words61[546-count_h];
          62 : wht <= words62[546-count_h];
          63 : wht <= words63[546-count_h];
          64 : wht <= words64[546-count_h];
          65 : wht <= words65[546-count_h];
          66 : wht <= words66[546-count_h];
          67 : wht <= words67[546-count_h];
          68 : wht <= words68[546-count_h];
          69 : wht <= words69[546-count_h];
          70 : wht <= words70[546-count_h];
          71 : wht <= words71[546-count_h];
          72 : wht <= words72[546-count_h];
          73 : wht <= words73[546-count_h];
          74 : wht <= words74[546-count_h];
          75 : wht <= words75[546-count_h];
          76 : wht <= words76[546-count_h];
          default: wht <= 1'b0;
        endcase
      end else begin
        wht <= 1'b0;
      end
    end
  end

  always @ (posedge clk) begin
    hs_out <= 1'b0;
    if (rst) begin
      count_h <= 10'b11_1111_1111;
      blank_h <= 1'b1;
    end else if (count_h < h_visible) begin
	  // horizontal visible
      count_h <= count_h + 1;
    end else if (count_h < h_frontporch) begin
	  // horizontal front porch
      count_h <= count_h + 1;
      blank_h <= 1'b1;
    end else if (count_h < h_sync) begin
	  // horizontal sync
      count_h <= count_h + 1;
	  hs_out <= 1'b1;
    end else if (count_h < h_backporch) begin
	  // horizontal back porch
      count_h <= count_h + 1;
    end else begin
      count_h <= 1;
      blank_h <= 1'b0;
    end
  end

  always @ (posedge clk) begin
    if (rst) begin
      count_v <= 15'b111_1111_1111_1111;
      blank_v <= 1'b1;
      vs_out  <= 1'b0;
    end else if (count_h >= h_backporch) begin
      if (count_v < v_visible) begin
        count_v <= count_v + 1;
      end else if (count_v < v_backporch) begin
        count_v <= count_v + 1;
        blank_v <= 1'b1;
        if (count_v > v_frontporch && count_v < v_sync) begin
          vs_out <= 1'b1;
        end else begin
          vs_out <= 1'b0;
        end
      end else begin
        count_v <= 1;
        blank_v <= 1'b0;
      end
    end
  end
  
endmodule
