
module vga(
	       input  clk,
	       input  rst,
	       output r0,
	       output r1,
	       output r2,
	       output r3,
	       output g0,
	       output g1,
	       output g2,
	       output g3,
	       output b0,
	       output b1,
	       output b2,
	       output b3,
	       output hs,
	       output vs
	       );

  localparam	  h_visible    = 640;
  localparam	  h_frontporch = 640 + 16;
  localparam	  h_sync       = 640 + 16 + 96;
  localparam	  h_backporch  = 640 + 16 + 96 + 47;

  // while h_sync is being sent, vertical counts h_sync pulses, for
  // porch and sync, it counts clocks
  localparam	  v_visible    = 480;
  localparam	  v_frontporch = 480 + 22;
  localparam	  v_sync       = 480 + 22 + 3;
  localparam	  v_backporch = 480 + 22 + 3 + 1;

  //   localparam smile001   = 59'b11111111111111111111111111111111111111111111111111111111111;
  //   localparam smile002   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile003   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile004   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile005   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile006   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile007   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile008   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile009   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile010   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile011   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile012   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile013   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile014   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile015   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile016   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile017   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile018   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile019   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile020   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile021   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile022   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile023   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile024   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile025   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile026   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile027   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile028   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile029   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile030   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile031   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile032   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile033   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile034   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile035   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile036   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile037   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile038   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile039   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile040   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile041   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile042   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile043   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile044   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile045   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile046   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile047   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile048   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile049   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile050   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile051   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile052   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile053   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile054   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile055   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile056   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile057   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile058   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile059   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile060   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile061   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile062   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile063   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile064   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile065   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile066   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile067   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile068   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile069   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile070   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile071   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile072   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile073   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile074   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile075   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile076   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile077   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile078   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile079   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile080   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile081   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile082   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile083   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile084   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile085   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile086   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile087   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile088   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile089   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile090   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile091   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile092   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile093   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile094   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile095   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile096   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile097   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile098   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile099   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile100   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile101   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile102   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile103   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile104   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile105   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile106   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile107   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile108   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile109   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile110   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile111   = 59'b10000000000000000000000000000000000000000000000000000000001;
  //   localparam smile112   = 59'b11111111111111111111111111111111111111111111111111111111111;
  localparam smile001  = 59'b00000000000000000000000000000000000000000000000000010000000;
  localparam smile002  = 59'b00000000000000000000000000000000000000000000000000111000000;
  localparam smile003  = 59'b00000000000000000000000000000000000000000000000000111110000;
  localparam smile004  = 59'b00000000000000000000000000000000000000000000000001111111000;
  localparam smile005  = 59'b00000000000000000000000000000000000000000000000011111111100;
  localparam smile006  = 59'b00000000000000000000000000000000000000000000000111111111110;
  localparam smile007  = 59'b00000000000000000000000000000000000000000000000111111111110;
  localparam smile008  = 59'b00000000000000000000000000000000000000000000001111111111100;
  localparam smile009  = 59'b00000000000000000000000000000000000000000000011111111111100;
  localparam smile010  = 59'b00000000000000000000000000000000000000000000011111111111000;
  localparam smile011  = 59'b00000000000000000000000000000000000000000000111111111110000;
  localparam smile012  = 59'b00000000000000000000000000000000000000000001111111111110000;
  localparam smile013  = 59'b00000000000000000000000000000000000000000001111111111100000;
  localparam smile014  = 59'b00000000000000000000000000000000000000000011111111111100000;
  localparam smile015  = 59'b00000000000000000000000000000000000000000011111111111000000;
  localparam smile016  = 59'b00000000000000000000000000000000000000000111111111110000000;
  localparam smile017  = 59'b00000000000000000000000000000000000000000111111111110000000;
  localparam smile018  = 59'b00000000000000000000000000000000000000001111111111100000000;
  localparam smile019  = 59'b00000000000000000000000000000000000000001111111111100000000;
  localparam smile020  = 59'b00000000000000000000000000000000000000011111111111000000000;
  localparam smile021  = 59'b00000000000000000000000000000000000000011111111111000000000;
  localparam smile022  = 59'b00000000000000000000000000000000000000111111111111000000000;
  localparam smile023  = 59'b00000000000000000000000000000000000000111111111110000000000;
  localparam smile024  = 59'b00000000000000000000000000000000000001111111111110000000000;
  localparam smile025  = 59'b00000000000000000000000000000000000001111111111100000000000;
  localparam smile026  = 59'b00000000000000000000000000000000000001111111111100000000000;
  localparam smile027  = 59'b00000000000000000000000000000000000011111111111100000000000;
  localparam smile028  = 59'b00000111111100000000000000000000000011111111111000000000000;
  localparam smile029  = 59'b00011111111111000000000000000000000011111111111000000000000;
  localparam smile030  = 59'b00111111111111100000000000000000000111111111111000000000000;
  localparam smile031  = 59'b01111111111111110000000000000000000111111111110000000000000;
  localparam smile032  = 59'b11111111111111111000000000000000000111111111110000000000000;
  localparam smile033  = 59'b11111111111111111000000000000000000111111111110000000000000;
  localparam smile034  = 59'b11111111111111111000000000000000001111111111110000000000000;
  localparam smile035  = 59'b11111111111111111100000000000000001111111111100000000000000;
  localparam smile036  = 59'b11111111111111111100000000000000001111111111100000000000000;
  localparam smile037  = 59'b11111111111111111100000000000000001111111111100000000000000;
  localparam smile038  = 59'b11111111111111111000000000000000001111111111100000000000000;
  localparam smile039  = 59'b11111111111111111000000000000000001111111111100000000000000;
  localparam smile040  = 59'b01111111111111111000000000000000011111111111000000000000000;
  localparam smile041  = 59'b01111111111111110000000000000000011111111111000000000000000;
  localparam smile042  = 59'b00111111111111100000000000000000011111111111000000000000000;
  localparam smile043  = 59'b00011111111111000000000000000000011111111111000000000000000;
  localparam smile044  = 59'b00000111111100000000000000000000011111111111000000000000000;
  localparam smile045  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile046  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile047  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile048  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile049  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile050  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile051  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile052  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile053  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile054  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile055  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile056  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile057  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile058  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile059  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile060  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile061  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile062  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile063  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile064  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile065  = 59'b00000000000000000000000000000000111111111110000000000000000;
  localparam smile066  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile067  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile068  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile069  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile070  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile071  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile072  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile073  = 59'b00000000000000000000000000000000011111111111000000000000000;
  localparam smile074  = 59'b00000000000000000000000000000000011111111111100000000000000;
  localparam smile075  = 59'b00000000000000000000000000000000001111111111100000000000000;
  localparam smile076  = 59'b00000000000000000000000000000000001111111111100000000000000;
  localparam smile077  = 59'b00000001110000000000000000000000001111111111100000000000000;
  localparam smile078  = 59'b00001111111110000000000000000000001111111111100000000000000;
  localparam smile079  = 59'b00011111111111100000000000000000001111111111110000000000000;
  localparam smile080  = 59'b00111111111111110000000000000000000111111111110000000000000;
  localparam smile081  = 59'b01111111111111110000000000000000000111111111110000000000000;
  localparam smile082  = 59'b11111111111111111000000000000000000111111111111000000000000;
  localparam smile083  = 59'b11111111111111111000000000000000000111111111111000000000000;
  localparam smile084  = 59'b11111111111111111000000000000000000011111111111000000000000;
  localparam smile085  = 59'b11111111111111111100000000000000000011111111111100000000000;
  localparam smile086  = 59'b11111111111111111100000000000000000011111111111100000000000;
  localparam smile087  = 59'b11111111111111111000000000000000000001111111111100000000000;
  localparam smile088  = 59'b11111111111111111000000000000000000001111111111110000000000;
  localparam smile089  = 59'b11111111111111111000000000000000000001111111111110000000000;
  localparam smile090  = 59'b01111111111111110000000000000000000000111111111110000000000;
  localparam smile091  = 59'b00111111111111110000000000000000000000111111111111000000000;
  localparam smile092  = 59'b00111111111111100000000000000000000000111111111111000000000;
  localparam smile093  = 59'b00001111111110000000000000000000000000011111111111100000000;
  localparam smile094  = 59'b00000011111000000000000000000000000000011111111111100000000;
  localparam smile095  = 59'b00000000000000000000000000000000000000001111111111110000000;
  localparam smile096  = 59'b00000000000000000000000000000000000000001111111111110000000;
  localparam smile097  = 59'b00000000000000000000000000000000000000000111111111111000000;
  localparam smile098  = 59'b00000000000000000000000000000000000000000111111111111000000;
  localparam smile099  = 59'b00000000000000000000000000000000000000000011111111111100000;
  localparam smile100  = 59'b00000000000000000000000000000000000000000001111111111110000;
  localparam smile101  = 59'b00000000000000000000000000000000000000000001111111111110000;
  localparam smile102  = 59'b00000000000000000000000000000000000000000000111111111111000;
  localparam smile103  = 59'b00000000000000000000000000000000000000000000111111111111000;
  localparam smile104  = 59'b00000000000000000000000000000000000000000000011111111111100;
  localparam smile105  = 59'b00000000000000000000000000000000000000000000001111111111110;
  localparam smile106  = 59'b00000000000000000000000000000000000000000000000111111111110;
  localparam smile107  = 59'b00000000000000000000000000000000000000000000000111111111111;
  localparam smile108  = 59'b00000000000000000000000000000000000000000000000011111111110;
  localparam smile109  = 59'b00000000000000000000000000000000000000000000000001111111100;
  localparam smile110  = 59'b00000000000000000000000000000000000000000000000000111111000;
  localparam smile111  = 59'b00000000000000000000000000000000000000000000000000011110000;
  localparam smile112  = 59'b00000000000000000000000000000000000000000000000000011000000;

  localparam words01  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000000000000000000000;
  localparam words02  = 588'b111100000000000111000000000000000000000000000000000000000000000000000000000000000111100000000000000111111111110000001110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000000000000;
  localparam words03  = 588'b011100000000001111000000000000000000000000000000000000000000000000000000000000000111110000000000001111111111110000001110000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words04  = 588'b011110000000011110000000000000000000000000000000000000000000000000000000000000001111110000000000011111100111110000001110000000011111110111111100000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words05  = 588'b001111000000011100000000000000000000000000000000000000000000000000000000000000001111111000000000111100000000010000001110000000111100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words06  = 588'b000111000000111100000000000000000000000000000000000000000000000000000000000000001110111000000000111000000000000000001110000001111000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words07  = 588'b000111100001111000001111110000000001100000000011000000110001111000000000000000011110111000000000111000000000000000001110000001110000000000000000000000000000110001111000001111111000000000110001111100000000000000000001100000011000111110000000111111111100000001111110000000000000000000001111111000000000000000000011000111110000000001100011110000001111110000000011110011111000000000111000000001111111000000001100011111000000111110000000000000000001100001111111111000000000000000000111111000000000111111000000000110000000001100000011100000000111110011110000011000111110000000001110001111111111;
  localparam words08  = 588'b000011110001110000111111111100000011110000000111100001111111111100000000000000011100111100000000111000000000000000001110000011110000000000000000000000000001111111111100111111111110000001111011111111000000000000000001110000111101111111100000111111111100000111111111100000000000000000111111111110000000000000000111111111111100000011111111111000111111111100000011111111111110000000111000000011111111100000011111111111100011111111000000000000000001110001111111111000000000000000011111111110000011111111110000001111000000011110000011100000011111111111110000111101111111100000001110001111111111;
  localparam words09  = 588'b000001110011110001111111111110000011110000000111100001111111111100000000000000111100011100000000111100000000000000001110000011110000000000000000000000000001111111111100111111111111000001111111111111100000000000000001110000111111111111110000111111111100001111111111110000000000000000111111111111000000000000000111111111111110000011111111111001111111111110000011111111111111000000111000000111111111110000011111111111110111111111100000000000000001110001111111111000000000000000111111111110000111111111111000001111000000011110000011100000111111111111110000111111111111110000001110001111111111;
  localparam words10  = 588'b000001111111100001111000001111000011110000000111100001111110000000000000000000111100011100000000111111000000000000001110000011100000000000000000000000000001111110000000100000001111000001111110000111100000000000000001110000111111000011110000011110000000001111000001111000000000000000100000001111000000000000000111111000011110000011111100000001111000001111000011111100001111000000111000001111000001111000011111100001111110000011100000000000000001110000111100000000000000000001111000000110000111100000111100001111000000011110000011100000111100001111110000111111000011110000001100000111100000;
  localparam words11  = 588'b000000111111000011110000001111000011110000000111100001111100000000000000000000111000011110000000011111111100000000001110000011100000000000000000000000000001111100000000000000000111100001111100000011100000000000000001110000111110000001110000011110000000011110000001111000000000000000000000000111100000000000000111110000001111000011111000000011110000001111000011111000000111100000111000011110000000111100011111000000111100000011110000000000000001110000111100000000000000000011110000000000001111000000111100001111000000011110000011100001111000000111110000111110000001110000000000000111100000;
  localparam words12  = 588'b000000011111000011100000000111100011110000000111100001111000000000000000000001111000001110000000001111111111100000001110000111100000000000000000000000000001111000000000000000000011100001111000000011110000000000000001110000111100000001111000011110000000011100000000111100000000000000000000000011100000000000000111100000000111000011110000000011100000000111100011110000000011100000111000011100000000011100011110000000111100000001110000000000000001110000111100000000000000000011100000000000001110000000011110001111000000011110000011100001110000000011110000111100000001111000000000000111100000;
  localparam words13  = 588'b000000011110000011100000000111100011110000000111100001111000000000000000000001110000001111000000000011111111110000001110000111100000000000000000000000000001111000000000000011111111100001111000000011110000000000000001110000111100000001111000011110000000011100000000111100000000000000000011111111100000000000000111100000000111000011110000000011100000000111100011110000000011100000111000011100000000011100011110000000111000000001110000000000000001110000111100000000000000000011100000000000001110000000011110001111000000011110000011100001110000000011110000111100000001111000000000000111100000;
  localparam words14  = 588'b000000011110000111100000000111100011110000000111100001111000000000000000000001110000001111000000000000001111111000001110000111100000000000000000000000000001111000000000011111111111100001111000000011110000000000000001110000111100000001111000011110000000111100000000111100000000000000011111111111100000000000000111100000000111100011110000000111100000000111100011110000000011110000111000111111111111111100011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000011110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words15  = 588'b000000011110000111100000000011100011110000000111100001111000000000000000000011110000000111000000000000000001111000001110000011100000000000000000000000000001111000000000111111111111100001111000000011110000000000000001110000111100000001111000011110000000111100000000011100000000000000111111111111100000000000000111100000000111100011110000000111100000000011100011110000000011110000111000111111111111111100011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000001110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words16  = 588'b000000011110000111100000000011100011110000000111100001111000000000000000000011111111111111100000000000000000111000001110000011110000000000000000000000000001111000000001111000000011100001111000000011110000000000000001110000111100000001111000011110000000111100000000011100000000000001111000000011100000000000000111100000000111100011110000000111100000000011100011110000000011110000111000111111111111111100011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000001110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words17  = 588'b000000011110000111100000000111100011110000000111100001111000000000000000000111111111111111100000000000000000111100001110000011110000000000000000000000000001111000000001110000000011100001111000000011110000000000000001110000111100000001111000011110000000111100000000111100000000000001110000000011100000000000000111100000000111100011110000000111100000000111100011110000000011110000111000111100000000000000011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000011110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words18  = 588'b000000011110000011100000000111100011110000000111100001111000000000000000000111111111111111100000000000000000111100001110000011110000000000000000000000000001111000000001110000000111100001111000000011110000000000000001110000111100000001111000001110000000011100000000111100000000000001110000000111100000000000000111100000000111000011110000000011100000000111100011110000000011100000111000011100000000000000011110000000111000000001110000000000000001110000011100000000000000000011100000000000001110000000011110001111000000011110000011100001110000000011110000111100000001111000000000000011100000;
  localparam words19  = 588'b000000011110000011110000000111000011110000000111100001111000000000000000000111000000000011110000000000000000111000001110000001111000000000000000000000000001111000000001110000000111100001111000000011110000000000000001110000111100000001111000001110000000011110000000111000000000000001110000000111100000000000000111100000000111000011110000000011110000000111000011110000000011100000111000011110000000000000011110000000111000000001110000000000000001110000011100000000000000000011110000000000001111000000011100001111000000011110000011100001110000000011110000111100000001111000000000000011100000;
  localparam words20  = 588'b000000011110000011110000001111000001110000001111100001111000000000000000001111000000000001110000110000000001111000001110000000111100000000011100000000000001111000000001110000001111100001111000000011110000000000000001110000111100000001111000001110000000011110000001111000000000000001110000001111100000000000000111110000001111000011110000000011110000001111000011111000000111100000111000011110000000000000011110000000111000000001110000000000000001110000011100000000000000000011110000000000001111000000111100000111000000111110000011100001111000000111110000111100000001111000000000000011100000;
  localparam words21  = 588'b000000011110000001111000011110000001111000011111100001111000000000000000001111000000000001111000111110000111111000001110000000111111100011111100000000000001111000000001111000011111100001111000000011110000000000000001110000111100000001111000001111111100001111000011110000000000000001111000011111100000000000000111111000011110000011110000000001111000011110000011111100001111000000111000001111100000111100011110000000111000000001110000000000000001110000011111111000000000000001111100001110000111100001111000000111100001111110000011100000111100001111110000111100000001111000000000000011111111;
  localparam words22  = 588'b000000011110000000111111111110000000111111111111100001111000000000000000001110000000000001111000111111111111110000001110000000011111111111111000000000000001111000000000111111111111100001111000000011110000000000000001110000111100000001111000001111111100000111111111110000000000000000111111111111100000000000000111111111111100000011110000000000111111111110000011111111111110000000111000000111111111111100011110000000111000000001110000000000000001110000011111111000000000000000111111111110000011111111111000000011111111111110000011100000011111111111110000111100000001111000000000000011111111;
  localparam words23  = 588'b000000011110000000011111111000000000011111110111100001111000000000000000011110000000000000111000011111111111100000001110000000000111111111110000000000000001111000000000011111110011100001111000000011110000000000000001110000111100000001111000000111111100000011111111000000000000000000011111110011100000000000000111101111111000000011110000000000011111111000000011110111111100000000111000000011111111111000011110000000111000000001110000000000000001110000001111111000000000000000011111111110000001111111100000000001111111011110000011100000001111111011110000111100000001111000000000000001111111;
  localparam words24  = 588'b000000000000000000000111100000000000000111000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000111110000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111000000000000000000000111100011100000000000000000000000000111100000000000000001110000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000011110000000000000011100000000000000000000000011100000000000000000000000000000000000000000000000;
  localparam words25  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words26  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words27  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words28  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words29  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words30  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words31  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words32  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words33  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words34  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words35  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words36  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words37  = 588'b001111001111100000000000111111100000000011000111110000000000001111100111100000111000000001111111000000000000000000001111111000000000110001111100000000000011111001111000000000000000110001111100000000000011111100000001110000000111000000011000000000000000110000111111111100000000000000110001111100000000000011111110000000000011111110000000000011111001111000000011111110000000000000001111111111000000011111100000000000000000001100011110000001111111000000000011111110000011111111110000001111111000000000110001111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words38  = 588'b001111011111111000000011111111111000000111101111111100000000111111111111100000111000000011111111100000000000000000111111111110000001111011111111000000001111111111111000000000000001111011111111000000001111111111000001110000001111000000111000000000000000111000111111111100000000000001111011111111000000000111111111000000000111111111000000001111111111111000001111111111100000000000001111111111000001111111111000000000000000011111111111000011111111100000001111111111100011111111110000111111111110000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words39  = 588'b001111111111111100000011111111111100000111111111111110000001111111111111100000111000000111111111110000000000000000111111111111000001111111111111100000011111111111111000000000000001111111111111100000011111111111100001111000001111100000111000000000000000111000111111111100000000000001111111111111100000001111111111100000001111111111100000011111111111111000011111111111100000000000001111111111000011111111111100000000000000011111111111000111111111110000011111111111100011111111110000111111111111000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words40  = 588'b001111110000111100000010000000111100000111111000011110000001111000011111100000111000001111000001111000000000000000100000001111000001111110000111100000011110000111111000000000000001111110000111100000011110000011110000111000001111100000111000000000000000111000011110000000000000000001111110000111100000011110000011110000011110000011110000011110000111111000011100000001000000000000000111100000000011110000011110000000000000011111100000001111000001111000011100000001000001111000000000100000001111000001111110000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words41  = 588'b001111100000011100000000000000011110000111110000001110000011110000001111100000111000011110000000111100000000000000000000000111100001111100000011100000111100000011111000000000000001111100000011100000111100000011110000111000011111100001111000000000000000111000011110000000000000000001111100000011100000111100000001111000111100000001111000111100000011111000011100000000000000000000000111100000000111100000011110000000000000011111000000011110000000111100011100000000000001111000000000000000000111100001111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words42  = 588'b001111000000011110000000000000001110000111100000001111000011100000000111100000111000011100000000011100000000000000000000000011100001111000000011110000111000000001111000000000000001111000000011110000111000000001111000111100011101100001110000000000000000111000011110000000000000000001111000000011110000111000000000111000111000000000111000111000000001111000111100000000000000000000000111100000000111000000001111000000000000011110000000011100000000011100111100000000000001111000000000000000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words43  = 588'b001111000000011110000000001111111110000111100000001111000011100000000111100000111000011100000000011100000000000000000011111111100001111000000011110000111000000001111000000000000001111000000011110000111000000001111000011100011101110001110000000000000000111000011110000000000000000001111000000011110000111000000000111000111000000000111000111000000001111000011110000000000000000000000111100000000111000000001111000000000000011110000000011100000000011100011110000000000001111000000000000011111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words44  = 588'b001111000000011110000001111111111110000111100000001111000111100000000111100000111000111111111111111100000000000000011111111111100001111000000011110001111000000001111000000000000001111000000011110001111000000001111000011100011101110011110000000000000000111000011110000000000000000001111000000011110001111111111111111001111111111111111001111000000001111000011111111000000000000000000111100000001111000000001111000000000000011110000000111111111111111100011111111000000001111000000000011111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words45  = 588'b001111000000011110000011111111111110000111100000001111000111100000000111100000111000111111111111111100000000000000111111111111100001111000000011110001111000000001111000000000000001111000000011110001111000000000111000011100111001110011100000000000000000111000011110000000000000000001111000000011110001111111111111111001111111111111111001111000000001111000001111111110000000000000000111100000001111000000000111000000000000011110000000111111111111111100001111111110000001111000000000111111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words46  = 588'b001111000000011110000111100000001110000111100000001111000111100000000111100000111000111111111111111100000000000001111000000011100001111000000011110001111000000001111000000000000001111000000011110001111000000000111000011110111000110011100000000000000000111000011110000000000000000001111000000011110001111111111111111001111111111111111001111000000001111000000011111111000000000000000111100000001111000000000111000000000000011110000000111111111111111100000011111111000001111000000001111000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words47  = 588'b001111000000011110000111000000001110000111100000001111000111100000000111100000111000111100000000000000000000000001110000000011100001111000000011110001111000000001111000000000000001111000000011110001111000000001111000001110111000111011100000000000000000111000011110000000000000000001111000000011110001111000000000000001111000000000000001111000000001111000000000001111100000000000000111100000001111000000001111000000000000011110000000111100000000000000000000001111100001111000000001110000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words48  = 588'b001111000000011110000111000000011110000111100000001111000011100000000111100000111000011100000000000000000000000001110000000111100001111000000011110000111000000001111000000000000001111000000011110000111000000001111000001110110000111111100000000000000000111000001110000000000000000001111000000011110000111000000000000000111000000000000000111000000001111000000000000011100000000000000011100000000111000000001111000000000000011110000000011100000000000000000000000011100000111000000001110000000111100001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words49  = 588'b001111000000011110000111000000011110000111100000001111000011100000000111100000111000011110000000000000000000000001110000000111100001111000000011110000111000000001111000000000000001111000000011110000111100000001110000001111110000111111000000000000000000111000001110000000000000000001111000000011110000111100000000000000111100000000000000111000000001111000000000000011100000000000000011100000000111100000001110000000000000011110000000011110000000000000000000000011100000111000000001110000000111100001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words50  = 588'b001111000000011110000111000000111110000111100000001111000011110000001111100000111000011110000000000000000000000001110000001111100001111000000011110000111100000011111000000000000001111000000011110000111100000011110000001111110000011111000000000000000000111000001110000000000000000001111000000011110000111100000000000000111100000000000000111100000011111000000000000011100000000000000011100000000111100000011110000000000000011110000000011110000000000000000000000011100000111000000001110000001111100001111000000000111000000000111000000000000000000000000000000000000000000000000000000000000000;
  localparam words51  = 588'b001111000000011110000111100001111110000111100000001111000001111000011111100000111000001111100000111100000000000001111000011111100001111000000011110000011110000111111000000000000001111000000011110000011110000111100000000111110000011111000000000000000000111000001111111100000000000001111000000011110000011111000001111000011111000001111000011110000111111000111100000111100000000000000011111111000011110000111100000000000000011110000000001111100000111100111100000111100000111111110001111000011111100001111000000000111111110000111100000000000000000000000000000000000000000000000000000000000000;
  localparam words52  = 588'b001111000000011110000011111111111110000111100000001111000000111111111111100000111000000111111111111100000000000000111111111111100001111000000011110000001111111111111000000000000001111000000011110000001111111111100000000111100000011111000000000000000000111000001111111100000000000001111000000011110000001111111111111000001111111111111000001111111111111000111111111111000000000000000011111111000001111111111100000000000000011110000000000111111111111100111111111111000000111111110000111111111111100001111000000000111111110000111100000000000000000000000000000000000000000000000000000000000000;
  localparam words53  = 588'b001111000000011110000001111111001110000111100000001111000000011111110111100000111000000011111111111000000000000000011111110011100001111000000011110000000111111101111000000000000001111000000011110000000111111110000000000111100000011110000000000000000000111000000111111100000000000001111000000011110000000111111111110000000111111111110000000111111101111000011111111110000000000000000001111111000000111111110000000000000000011110000000000011111111111000011111111110000000011111110000011111110011100001111000000000011111110000111100000000000000000000000000000000000000000000000000000000000000;
  localparam words54  = 588'b000000000000000000000000011100000000000000000000000000000000000111000000000000000000000000011111000000000000000000000111000000000000000000000000000000000001110000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000111110000000000001110000000000000011111000000000000000000000000000000000001111000000000000000000000000000000000000011111000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  wire            blank;
  reg             blank_h;
  reg             blank_v;

  assign blank = (blank_h | blank_v);

  // 2^10  = 1024
  reg [9:0]       count_h;
  // 2^15 = 32768
  reg [14:0]      count_v;

  

  reg             red;
  reg             grn;
  wire            blu;
  wire            wht;
  reg             hs_out;
  reg             vs_out;

  reg [3:0]       fb[3:0];

  reg [53:0]     row;

  assign r0 = red;
  assign r1 = red;
  assign r2 = red;
  assign r3 = red;
  assign b0 = blu;
  assign b1 = blu;
  assign b2 = blu;
  assign b3 = blu;
  assign g0 = grn;
  assign g1 = grn;
  assign g2 = grn;
  assign g3 = grn;
  assign hs = !hs_out;
  assign vs = !vs_out;

  always @ (posedge clk) begin
    if (rst) begin
      red <= 1'b0;
      grn <= 1'b0;
    end else begin
      red <= wht;
      grn <= wht;
    end
  end

  //   assign red = wht;
  //   assign grn = wht;

  assign blu = (blank) ? 1'b0 : 1'b1;

  assign wht            = (count_h < 20 || count_h > 607) ? 1'b0 :
//                           (count_v == 100 && count_h < 79) ? smile001[78-count_h] :
//                           (count_v == 101 && count_h < 79) ? smile002[78-count_h] :
//                           (count_v == 102 && count_h < 79) ? smile003[78-count_h] :
//                           (count_v == 103 && count_h < 79) ? smile004[78-count_h] :
//                           (count_v == 104 && count_h < 79) ? smile005[78-count_h] :
//                           (count_v == 105 && count_h < 79) ? smile006[78-count_h] :
//                           (count_v == 106 && count_h < 79) ? smile007[78-count_h] :
//                           (count_v == 107 && count_h < 79) ? smile008[78-count_h] :
//                           (count_v == 108 && count_h < 79) ? smile009[78-count_h] :
//                           (count_v == 109 && count_h < 79) ? smile010[78-count_h] :
//                           (count_v == 110 && count_h < 79) ? smile011[78-count_h] :
//                           (count_v == 111 && count_h < 79) ? smile012[78-count_h] :
//                           (count_v == 112 && count_h < 79) ? smile013[78-count_h] :
//                           (count_v == 113 && count_h < 79) ? smile014[78-count_h] :
//                           (count_v == 114 && count_h < 79) ? smile015[78-count_h] :
//                           (count_v == 115 && count_h < 79) ? smile016[78-count_h] :
//                           (count_v == 116 && count_h < 79) ? smile017[78-count_h] :
//                           (count_v == 117 && count_h < 79) ? smile018[78-count_h] :
//                           (count_v == 118 && count_h < 79) ? smile019[78-count_h] :
//                           (count_v == 119 && count_h < 79) ? smile020[78-count_h] :
//                           (count_v == 120 && count_h < 79) ? smile021[78-count_h] :
//                           (count_v == 121 && count_h < 79) ? smile022[78-count_h] :
//                           (count_v == 122 && count_h < 79) ? smile023[78-count_h] :
//                           (count_v == 123 && count_h < 79) ? smile024[78-count_h] :
//                           (count_v == 124 && count_h < 79) ? smile025[78-count_h] :
//                           (count_v == 125 && count_h < 79) ? smile026[78-count_h] :
//                           (count_v == 126 && count_h < 79) ? smile027[78-count_h] :
//                           (count_v == 127 && count_h < 79) ? smile028[78-count_h] :
//                           (count_v == 128 && count_h < 79) ? smile029[78-count_h] :
//                           (count_v == 129 && count_h < 79) ? smile030[78-count_h] :
//                           (count_v == 130 && count_h < 79) ? smile031[78-count_h] :
//                           (count_v == 131 && count_h < 79) ? smile032[78-count_h] :
//                           (count_v == 132 && count_h < 79) ? smile033[78-count_h] :
//                           (count_v == 133 && count_h < 79) ? smile034[78-count_h] :
//                           (count_v == 134 && count_h < 79) ? smile035[78-count_h] :
//                           (count_v == 135 && count_h < 79) ? smile036[78-count_h] :
//                           (count_v == 136 && count_h < 79) ? smile037[78-count_h] :
//                           (count_v == 137 && count_h < 79) ? smile038[78-count_h] :
//                           (count_v == 138 && count_h < 79) ? smile039[78-count_h] :
//                           (count_v == 139 && count_h < 79) ? smile040[78-count_h] :
//                           (count_v == 140 && count_h < 79) ? smile041[78-count_h] :
//                           (count_v == 141 && count_h < 79) ? smile042[78-count_h] :
//                           (count_v == 142 && count_h < 79) ? smile043[78-count_h] :
//                           (count_v == 143 && count_h < 79) ? smile044[78-count_h] :
//                           (count_v == 144 && count_h < 79) ? smile045[78-count_h] :
//                           (count_v == 145 && count_h < 79) ? smile046[78-count_h] :
//                           (count_v == 146 && count_h < 79) ? smile047[78-count_h] :
//                           (count_v == 147 && count_h < 79) ? smile048[78-count_h] :
//                           (count_v == 148 && count_h < 79) ? smile049[78-count_h] :
//                           (count_v == 149 && count_h < 79) ? smile050[78-count_h] :
//                           (count_v == 150 && count_h < 79) ? smile051[78-count_h] :
//                           (count_v == 151 && count_h < 79) ? smile052[78-count_h] :
//                           (count_v == 152 && count_h < 79) ? smile053[78-count_h] :
//                           (count_v == 153 && count_h < 79) ? smile054[78-count_h] :
//                           (count_v == 154 && count_h < 79) ? smile055[78-count_h] :
//                           (count_v == 155 && count_h < 79) ? smile056[78-count_h] :
//                           (count_v == 156 && count_h < 79) ? smile057[78-count_h] :
//                           (count_v == 157 && count_h < 79) ? smile058[78-count_h] :
//                           (count_v == 158 && count_h < 79) ? smile059[78-count_h] :
//                           (count_v == 159 && count_h < 79) ? smile060[78-count_h] :
//                           (count_v == 160 && count_h < 79) ? smile061[78-count_h] :
//                           (count_v == 161 && count_h < 79) ? smile062[78-count_h] :
//                           (count_v == 162 && count_h < 79) ? smile063[78-count_h] :
//                           (count_v == 163 && count_h < 79) ? smile064[78-count_h] :
//                           (count_v == 164 && count_h < 79) ? smile065[78-count_h] :
//                           (count_v == 165 && count_h < 79) ? smile066[78-count_h] :
//                           (count_v == 166 && count_h < 79) ? smile067[78-count_h] :
//                           (count_v == 167 && count_h < 79) ? smile068[78-count_h] :
//                           (count_v == 168 && count_h < 79) ? smile069[78-count_h] :
//                           (count_v == 169 && count_h < 79) ? smile070[78-count_h] :
//                           (count_v == 170 && count_h < 79) ? smile071[78-count_h] :
//                           (count_v == 171 && count_h < 79) ? smile072[78-count_h] :
//                           (count_v == 172 && count_h < 79) ? smile073[78-count_h] :
//                           (count_v == 173 && count_h < 79) ? smile074[78-count_h] :
//                           (count_v == 174 && count_h < 79) ? smile075[78-count_h] :
//                           (count_v == 175 && count_h < 79) ? smile076[78-count_h] :
//                           (count_v == 176 && count_h < 79) ? smile077[78-count_h] :
//                           (count_v == 177 && count_h < 79) ? smile078[78-count_h] :
//                           (count_v == 178 && count_h < 79) ? smile079[78-count_h] :
//                           (count_v == 179 && count_h < 79) ? smile080[78-count_h] :
//                           (count_v == 180 && count_h < 79) ? smile081[78-count_h] :
//                           (count_v == 181 && count_h < 79) ? smile082[78-count_h] :
//                           (count_v == 182 && count_h < 79) ? smile083[78-count_h] :
//                           (count_v == 183 && count_h < 79) ? smile084[78-count_h] :
//                           (count_v == 184 && count_h < 79) ? smile085[78-count_h] :
//                           (count_v == 185 && count_h < 79) ? smile086[78-count_h] :
//                           (count_v == 186 && count_h < 79) ? smile087[78-count_h] :
//                           (count_v == 187 && count_h < 79) ? smile088[78-count_h] :
//                           (count_v == 188 && count_h < 79) ? smile089[78-count_h] :
//                           (count_v == 189 && count_h < 79) ? smile090[78-count_h] :
//                           (count_v == 190 && count_h < 79) ? smile091[78-count_h] :
//                           (count_v == 191 && count_h < 79) ? smile092[78-count_h] :
//                           (count_v == 192 && count_h < 79) ? smile093[78-count_h] :
//                           (count_v == 193 && count_h < 79) ? smile094[78-count_h] :
//                           (count_v == 194 && count_h < 79) ? smile095[78-count_h] :
//                           (count_v == 195 && count_h < 79) ? smile096[78-count_h] :
//                           (count_v == 196 && count_h < 79) ? smile097[78-count_h] :
//                           (count_v == 197 && count_h < 79) ? smile098[78-count_h] :
//                           (count_v == 198 && count_h < 79) ? smile099[78-count_h] :
//                           (count_v == 199 && count_h < 79) ? smile100[78-count_h] :
//                           (count_v == 200 && count_h < 79) ? smile101[78-count_h] :
//                           (count_v == 201 && count_h < 79) ? smile102[78-count_h] :
//                           (count_v == 202 && count_h < 79) ? smile103[78-count_h] :
//                           (count_v == 203 && count_h < 79) ? smile104[78-count_h] :
//                           (count_v == 204 && count_h < 79) ? smile105[78-count_h] :
//                           (count_v == 205 && count_h < 79) ? smile106[78-count_h] :
//                           (count_v == 206 && count_h < 79) ? smile107[78-count_h] :
//                           (count_v == 207 && count_h < 79) ? smile108[78-count_h] :
//                           (count_v == 208 && count_h < 79) ? smile109[78-count_h] :
//                           (count_v == 209 && count_h < 79) ? smile110[78-count_h] :
//                           (count_v == 210 && count_h < 79) ? smile111[78-count_h] :
//                           (count_v == 211 && count_h < 79) ? smile112[78-count_h] :
                          (row[0] == 1'b1) ? words01[607-count_h] :
                          (row[1] == 1'b1) ? words02[607-count_h] :
                          (row[2] == 1'b1) ? words03[607-count_h] :
                          (row[3] == 1'b1) ? words04[607-count_h] :
                          (row[4] == 1'b1) ? words05[607-count_h] :
                          (row[5] == 1'b1) ? words06[607-count_h] :
                          (row[6] == 1'b1) ? words07[607-count_h] :
                          (row[7] == 1'b1) ? words08[607-count_h] :
                          (row[8] == 1'b1) ? words09[607-count_h] :
                          (row[9] == 1'b1) ? words10[607-count_h] :
                          (row[10] == 1'b1) ? words11[607-count_h] :
                          (row[11] == 1'b1) ? words12[607-count_h] :
                          (row[12] == 1'b1) ? words13[607-count_h] :
                          (row[13] == 1'b1) ? words14[607-count_h] :
                          (row[14] == 1'b1) ? words15[607-count_h] :
                          (row[15] == 1'b1) ? words16[607-count_h] :
                          (row[16] == 1'b1) ? words17[607-count_h] :
                          (row[17] == 1'b1) ? words18[607-count_h] :
                          (row[18] == 1'b1) ? words19[607-count_h] :
                          (row[19] == 1'b1) ? words20[607-count_h] :
                          (row[20] == 1'b1) ? words21[607-count_h] :
                          (row[21] == 1'b1) ? words22[607-count_h] :
                          (row[22] == 1'b1) ? words23[607-count_h] :
                          (row[23] == 1'b1) ? words24[607-count_h] :
                          (row[24] == 1'b1) ? words25[607-count_h] :
                          (row[25] == 1'b1) ? words26[607-count_h] :
                          (row[26] == 1'b1) ? words27[607-count_h] :
                          (row[27] == 1'b1) ? words28[607-count_h] :
                          (row[28] == 1'b1) ? words29[607-count_h] :
                          (row[29] == 1'b1) ? words30[607-count_h] :
                          (row[30] == 1'b1) ? words31[607-count_h] :
                          (row[31] == 1'b1) ? words32[607-count_h] :
                          (row[32] == 1'b1) ? words33[607-count_h] :
                          (row[33] == 1'b1) ? words34[607-count_h] :
                          (row[34] == 1'b1) ? words35[607-count_h] :
                          (row[35] == 1'b1) ? words36[607-count_h] :
                          (row[36] == 1'b1) ? words37[607-count_h] :
                          (row[37] == 1'b1) ? words38[607-count_h] :
                          (row[38] == 1'b1) ? words39[607-count_h] :
                          (row[39] == 1'b1) ? words40[607-count_h] :
                          (row[40] == 1'b1) ? words41[607-count_h] :
                          (row[41] == 1'b1) ? words42[607-count_h] :
                          (row[42] == 1'b1) ? words43[607-count_h] :
                          (row[43] == 1'b1) ? words44[607-count_h] :
                          (row[44] == 1'b1) ? words45[607-count_h] :
                          (row[45] == 1'b1) ? words46[607-count_h] :
                          (row[46] == 1'b1) ? words47[607-count_h] :
                          (row[47] == 1'b1) ? words48[607-count_h] :
                          (row[48] == 1'b1) ? words49[607-count_h] :
                          (row[49] == 1'b1) ? words50[607-count_h] :
                          (row[50] == 1'b1) ? words51[607-count_h] :
                          (row[51] == 1'b1) ? words52[607-count_h] :
                          (row[52] == 1'b1) ? words53[607-count_h] :
                          (row[53] == 1'b1) ? words54[607-count_h] :
                          1'b0;

  always @ (posedge clk) begin
    hs_out <= 1'b0;
    if (rst) begin
      count_h <= 10'b11_1111_1111;
      blank_h <= 1'b1;
    end else if (count_h < h_visible) begin
	  // horizontal visible
      count_h <= count_h + 1;
    end else if (count_h < h_frontporch) begin
	  // horizontal front porch
      count_h <= count_h + 1;
      blank_h <= 1'b1;
    end else if (count_h < h_sync) begin
	  // horizontal sync
      count_h <= count_h + 1;
	  hs_out <= 1'b1;
    end else if (count_h < h_backporch) begin
	  // horizontal back porch
      count_h <= count_h + 1;
    end else begin
      count_h <= 1;
      blank_h <= 1'b0;
    end
  end

  always @ (posedge clk) begin
    if (rst) begin
      count_v              <= 15'b111_1111_1111_1111;
      blank_v              <= 1'b1;
      vs_out               <= 1'b0;
      row                  <= 0;
      end else if (count_h >= h_backporch) begin
      if (count_v < v_visible) begin
        count_v <= count_v + 1;
        if (count_v > 299 && count_v < 354) begin
          row    <= row << 1;
          row[0] <= 1'b0;
        end else begin
          row[0] <= 1'b1;
        end
      end else if (count_v < v_backporch) begin
        count_v <= count_v + 1;
        blank_v <= 1'b1;
        if (count_v > v_frontporch && count_v < v_sync) begin
          vs_out <= 1'b1;
        end else begin
          vs_out <= 1'b0;
        end
      end else begin
        count_v <= 1;
        blank_v <= 1'b0;
      end
    end
  end
  
endmodule
