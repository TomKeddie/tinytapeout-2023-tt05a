module vga(
	       input  clk,
	       input  rst,
	       output r0,
	       output r1,
	       output r2,
	       output r3,
	       output g0,
	       output g1,
	       output g2,
	       output g3,
	       output b0,
	       output b1,
	       output b2,
	       output b3,
	       output hs,
	       output vs
	       );

  localparam	  h_visible    = 640;
  localparam	  h_frontporch = 640 + 16;
  localparam	  h_sync       = 640 + 16 + 96;
  localparam	  h_backporch  = 640 + 16 + 96 + 47;

  // while h_sync is being sent, vertical counts h_sync pulses, for
  // porch and sync, it counts clocks
  localparam	  v_visible    = 480;
  localparam	  v_frontporch = 480 + 22;
  localparam	  v_sync       = 480 + 22 + 3;
  localparam	  v_backporch = 480 + 22 + 3 + 1;

  localparam smile001   = 59'b11111111111111111111111111111111111111111111111111111111111;
  localparam smile002   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile003   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile004   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile005   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile006   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile007   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile008   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile009   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile010   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile011   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile012   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile013   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile014   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile015   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile016   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile017   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile018   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile019   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile020   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile021   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile022   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile023   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile024   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile025   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile026   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile027   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile028   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile029   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile030   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile031   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile032   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile033   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile034   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile035   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile036   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile037   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile038   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile039   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile040   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile041   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile042   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile043   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile044   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile045   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile046   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile047   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile048   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile049   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile050   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile051   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile052   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile053   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile054   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile055   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile056   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile057   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile058   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile059   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile060   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile061   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile062   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile063   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile064   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile065   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile066   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile067   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile068   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile069   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile070   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile071   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile072   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile073   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile074   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile075   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile076   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile077   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile078   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile079   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile080   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile081   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile082   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile083   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile084   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile085   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile086   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile087   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile088   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile089   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile090   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile091   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile092   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile093   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile094   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile095   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile096   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile097   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile098   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile099   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile100   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile101   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile102   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile103   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile104   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile105   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile106   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile107   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile108   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile109   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile110   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile111   = 59'b10000000000000000000000000000000000000000000000000000000001;
  localparam smile112   = 59'b11111111111111111111111111111111111111111111111111111111111;
  // localparam smile001  = 59'b00000000000000000000000000000000000000000000000000010000000;
  // localparam smile002  = 59'b00000000000000000000000000000000000000000000000000111000000;
  // localparam smile003  = 59'b00000000000000000000000000000000000000000000000000111110000;
  // localparam smile004  = 59'b00000000000000000000000000000000000000000000000001111111000;
  // localparam smile005  = 59'b00000000000000000000000000000000000000000000000011111111100;
  // localparam smile006  = 59'b00000000000000000000000000000000000000000000000111111111110;
  // localparam smile007  = 59'b00000000000000000000000000000000000000000000000111111111110;
  // localparam smile008  = 59'b00000000000000000000000000000000000000000000001111111111100;
  // localparam smile009  = 59'b00000000000000000000000000000000000000000000011111111111100;
  // localparam smile010  = 59'b00000000000000000000000000000000000000000000011111111111000;
  // localparam smile011  = 59'b00000000000000000000000000000000000000000000111111111110000;
  // localparam smile012  = 59'b00000000000000000000000000000000000000000001111111111110000;
  // localparam smile013  = 59'b00000000000000000000000000000000000000000001111111111100000;
  // localparam smile014  = 59'b00000000000000000000000000000000000000000011111111111100000;
  // localparam smile015  = 59'b00000000000000000000000000000000000000000011111111111000000;
  // localparam smile016  = 59'b00000000000000000000000000000000000000000111111111110000000;
  // localparam smile017  = 59'b00000000000000000000000000000000000000000111111111110000000;
  // localparam smile018  = 59'b00000000000000000000000000000000000000001111111111100000000;
  // localparam smile019  = 59'b00000000000000000000000000000000000000001111111111100000000;
  // localparam smile020  = 59'b00000000000000000000000000000000000000011111111111000000000;
  // localparam smile021  = 59'b00000000000000000000000000000000000000011111111111000000000;
  // localparam smile022  = 59'b00000000000000000000000000000000000000111111111111000000000;
  // localparam smile023  = 59'b00000000000000000000000000000000000000111111111110000000000;
  // localparam smile024  = 59'b00000000000000000000000000000000000001111111111110000000000;
  // localparam smile025  = 59'b00000000000000000000000000000000000001111111111100000000000;
  // localparam smile026  = 59'b00000000000000000000000000000000000001111111111100000000000;
  // localparam smile027  = 59'b00000000000000000000000000000000000011111111111100000000000;
  // localparam smile028  = 59'b00000111111100000000000000000000000011111111111000000000000;
  // localparam smile029  = 59'b00011111111111000000000000000000000011111111111000000000000;
  // localparam smile030  = 59'b00111111111111100000000000000000000111111111111000000000000;
  // localparam smile031  = 59'b01111111111111110000000000000000000111111111110000000000000;
  // localparam smile032  = 59'b11111111111111111000000000000000000111111111110000000000000;
  // localparam smile033  = 59'b11111111111111111000000000000000000111111111110000000000000;
  // localparam smile034  = 59'b11111111111111111000000000000000001111111111110000000000000;
  // localparam smile035  = 59'b11111111111111111100000000000000001111111111100000000000000;
  // localparam smile036  = 59'b11111111111111111100000000000000001111111111100000000000000;
  // localparam smile037  = 59'b11111111111111111100000000000000001111111111100000000000000;
  // localparam smile038  = 59'b11111111111111111000000000000000001111111111100000000000000;
  // localparam smile039  = 59'b11111111111111111000000000000000001111111111100000000000000;
  // localparam smile040  = 59'b01111111111111111000000000000000011111111111000000000000000;
  // localparam smile041  = 59'b01111111111111110000000000000000011111111111000000000000000;
  // localparam smile042  = 59'b00111111111111100000000000000000011111111111000000000000000;
  // localparam smile043  = 59'b00011111111111000000000000000000011111111111000000000000000;
  // localparam smile044  = 59'b00000111111100000000000000000000011111111111000000000000000;
  // localparam smile045  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile046  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile047  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile048  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile049  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile050  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile051  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile052  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile053  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile054  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile055  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile056  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile057  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile058  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile059  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile060  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile061  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile062  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile063  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile064  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile065  = 59'b00000000000000000000000000000000111111111110000000000000000;
  // localparam smile066  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile067  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile068  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile069  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile070  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile071  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile072  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile073  = 59'b00000000000000000000000000000000011111111111000000000000000;
  // localparam smile074  = 59'b00000000000000000000000000000000011111111111100000000000000;
  // localparam smile075  = 59'b00000000000000000000000000000000001111111111100000000000000;
  // localparam smile076  = 59'b00000000000000000000000000000000001111111111100000000000000;
  // localparam smile077  = 59'b00000001110000000000000000000000001111111111100000000000000;
  // localparam smile078  = 59'b00001111111110000000000000000000001111111111100000000000000;
  // localparam smile079  = 59'b00011111111111100000000000000000001111111111110000000000000;
  // localparam smile080  = 59'b00111111111111110000000000000000000111111111110000000000000;
  // localparam smile081  = 59'b01111111111111110000000000000000000111111111110000000000000;
  // localparam smile082  = 59'b11111111111111111000000000000000000111111111111000000000000;
  // localparam smile083  = 59'b11111111111111111000000000000000000111111111111000000000000;
  // localparam smile084  = 59'b11111111111111111000000000000000000011111111111000000000000;
  // localparam smile085  = 59'b11111111111111111100000000000000000011111111111100000000000;
  // localparam smile086  = 59'b11111111111111111100000000000000000011111111111100000000000;
  // localparam smile087  = 59'b11111111111111111000000000000000000001111111111100000000000;
  // localparam smile088  = 59'b11111111111111111000000000000000000001111111111110000000000;
  // localparam smile089  = 59'b11111111111111111000000000000000000001111111111110000000000;
  // localparam smile090  = 59'b01111111111111110000000000000000000000111111111110000000000;
  // localparam smile091  = 59'b00111111111111110000000000000000000000111111111111000000000;
  // localparam smile092  = 59'b00111111111111100000000000000000000000111111111111000000000;
  // localparam smile093  = 59'b00001111111110000000000000000000000000011111111111100000000;
  // localparam smile094  = 59'b00000011111000000000000000000000000000011111111111100000000;
  // localparam smile095  = 59'b00000000000000000000000000000000000000001111111111110000000;
  // localparam smile096  = 59'b00000000000000000000000000000000000000001111111111110000000;
  // localparam smile097  = 59'b00000000000000000000000000000000000000000111111111111000000;
  // localparam smile098  = 59'b00000000000000000000000000000000000000000111111111111000000;
  // localparam smile099  = 59'b00000000000000000000000000000000000000000011111111111100000;
  // localparam smile100  = 59'b00000000000000000000000000000000000000000001111111111110000;
  // localparam smile101  = 59'b00000000000000000000000000000000000000000001111111111110000;
  // localparam smile102  = 59'b00000000000000000000000000000000000000000000111111111111000;
  // localparam smile103  = 59'b00000000000000000000000000000000000000000000111111111111000;
  // localparam smile104  = 59'b00000000000000000000000000000000000000000000011111111111100;
  // localparam smile105  = 59'b00000000000000000000000000000000000000000000001111111111110;
  // localparam smile106  = 59'b00000000000000000000000000000000000000000000000111111111110;
  // localparam smile107  = 59'b00000000000000000000000000000000000000000000000111111111111;
  // localparam smile108  = 59'b00000000000000000000000000000000000000000000000011111111110;
  // localparam smile109  = 59'b00000000000000000000000000000000000000000000000001111111100;
  // localparam smile110  = 59'b00000000000000000000000000000000000000000000000000111111000;
  // localparam smile111  = 59'b00000000000000000000000000000000000000000000000000011110000;
  // localparam smile112  = 59'b00000000000000000000000000000000000000000000000000011000000;

  localparam words01  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000000000000000000000;
  localparam words02  = 588'b111100000000000111000000000000000000000000000000000000000000000000000000000000000111100000000000000111111111110000001110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000000000000;
  localparam words03  = 588'b011100000000001111000000000000000000000000000000000000000000000000000000000000000111110000000000001111111111110000001110000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words04  = 588'b011110000000011110000000000000000000000000000000000000000000000000000000000000001111110000000000011111100111110000001110000000011111110111111100000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000001110000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words05  = 588'b001111000000011100000000000000000000000000000000000000000000000000000000000000001111111000000000111100000000010000001110000000111100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words06  = 588'b000111000000111100000000000000000000000000000000000000000000000000000000000000001110111000000000111000000000000000001110000001111000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000000000000000001110000111100000;
  localparam words07  = 588'b000111100001111000001111110000000001100000000011000000110001111000000000000000011110111000000000111000000000000000001110000001110000000000000000000000000000110001111000001111111000000000110001111100000000000000000001100000011000111110000000111111111100000001111110000000000000000000001111111000000000000000000011000111110000000001100011110000001111110000000011110011111000000000111000000001111111000000001100011111000000111110000000000000000001100001111111111000000000000000000111111000000000111111000000000110000000001100000011100000000111110011110000011000111110000000001110001111111111;
  localparam words08  = 588'b000011110001110000111111111100000011110000000111100001111111111100000000000000011100111100000000111000000000000000001110000011110000000000000000000000000001111111111100111111111110000001111011111111000000000000000001110000111101111111100000111111111100000111111111100000000000000000111111111110000000000000000111111111111100000011111111111000111111111100000011111111111110000000111000000011111111100000011111111111100011111111000000000000000001110001111111111000000000000000011111111110000011111111110000001111000000011110000011100000011111111111110000111101111111100000001110001111111111;
  localparam words09  = 588'b000001110011110001111111111110000011110000000111100001111111111100000000000000111100011100000000111100000000000000001110000011110000000000000000000000000001111111111100111111111111000001111111111111100000000000000001110000111111111111110000111111111100001111111111110000000000000000111111111111000000000000000111111111111110000011111111111001111111111110000011111111111111000000111000000111111111110000011111111111110111111111100000000000000001110001111111111000000000000000111111111110000111111111111000001111000000011110000011100000111111111111110000111111111111110000001110001111111111;
  localparam words10  = 588'b000001111111100001111000001111000011110000000111100001111110000000000000000000111100011100000000111111000000000000001110000011100000000000000000000000000001111110000000100000001111000001111110000111100000000000000001110000111111000011110000011110000000001111000001111000000000000000100000001111000000000000000111111000011110000011111100000001111000001111000011111100001111000000111000001111000001111000011111100001111110000011100000000000000001110000111100000000000000000001111000000110000111100000111100001111000000011110000011100000111100001111110000111111000011110000001100000111100000;
  localparam words11  = 588'b000000111111000011110000001111000011110000000111100001111100000000000000000000111000011110000000011111111100000000001110000011100000000000000000000000000001111100000000000000000111100001111100000011100000000000000001110000111110000001110000011110000000011110000001111000000000000000000000000111100000000000000111110000001111000011111000000011110000001111000011111000000111100000111000011110000000111100011111000000111100000011110000000000000001110000111100000000000000000011110000000000001111000000111100001111000000011110000011100001111000000111110000111110000001110000000000000111100000;
  localparam words12  = 588'b000000011111000011100000000111100011110000000111100001111000000000000000000001111000001110000000001111111111100000001110000111100000000000000000000000000001111000000000000000000011100001111000000011110000000000000001110000111100000001111000011110000000011100000000111100000000000000000000000011100000000000000111100000000111000011110000000011100000000111100011110000000011100000111000011100000000011100011110000000111100000001110000000000000001110000111100000000000000000011100000000000001110000000011110001111000000011110000011100001110000000011110000111100000001111000000000000111100000;
  localparam words13  = 588'b000000011110000011100000000111100011110000000111100001111000000000000000000001110000001111000000000011111111110000001110000111100000000000000000000000000001111000000000000011111111100001111000000011110000000000000001110000111100000001111000011110000000011100000000111100000000000000000011111111100000000000000111100000000111000011110000000011100000000111100011110000000011100000111000011100000000011100011110000000111000000001110000000000000001110000111100000000000000000011100000000000001110000000011110001111000000011110000011100001110000000011110000111100000001111000000000000111100000;
  localparam words14  = 588'b000000011110000111100000000111100011110000000111100001111000000000000000000001110000001111000000000000001111111000001110000111100000000000000000000000000001111000000000011111111111100001111000000011110000000000000001110000111100000001111000011110000000111100000000111100000000000000011111111111100000000000000111100000000111100011110000000111100000000111100011110000000011110000111000111111111111111100011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000011110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words15  = 588'b000000011110000111100000000011100011110000000111100001111000000000000000000011110000000111000000000000000001111000001110000011100000000000000000000000000001111000000000111111111111100001111000000011110000000000000001110000111100000001111000011110000000111100000000011100000000000000111111111111100000000000000111100000000111100011110000000111100000000011100011110000000011110000111000111111111111111100011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000001110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words16  = 588'b000000011110000111100000000011100011110000000111100001111000000000000000000011111111111111100000000000000000111000001110000011110000000000000000000000000001111000000001111000000011100001111000000011110000000000000001110000111100000001111000011110000000111100000000011100000000000001111000000011100000000000000111100000000111100011110000000111100000000011100011110000000011110000111000111111111111111100011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000001110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words17  = 588'b000000011110000111100000000111100011110000000111100001111000000000000000000111111111111111100000000000000000111100001110000011110000000000000000000000000001111000000001110000000011100001111000000011110000000000000001110000111100000001111000011110000000111100000000111100000000000001110000000011100000000000000111100000000111100011110000000111100000000111100011110000000011110000111000111100000000000000011110000000111000000001110000000000000001110000111100000000000000000111100000000000011110000000011110001111000000011110000011100011110000000011110000111100000001111000000000000111100000;
  localparam words18  = 588'b000000011110000011100000000111100011110000000111100001111000000000000000000111111111111111100000000000000000111100001110000011110000000000000000000000000001111000000001110000000111100001111000000011110000000000000001110000111100000001111000001110000000011100000000111100000000000001110000000111100000000000000111100000000111000011110000000011100000000111100011110000000011100000111000011100000000000000011110000000111000000001110000000000000001110000011100000000000000000011100000000000001110000000011110001111000000011110000011100001110000000011110000111100000001111000000000000011100000;
  localparam words19  = 588'b000000011110000011110000000111000011110000000111100001111000000000000000000111000000000011110000000000000000111000001110000001111000000000000000000000000001111000000001110000000111100001111000000011110000000000000001110000111100000001111000001110000000011110000000111000000000000001110000000111100000000000000111100000000111000011110000000011110000000111000011110000000011100000111000011110000000000000011110000000111000000001110000000000000001110000011100000000000000000011110000000000001111000000011100001111000000011110000011100001110000000011110000111100000001111000000000000011100000;
  localparam words20  = 588'b000000011110000011110000001111000001110000001111100001111000000000000000001111000000000001110000110000000001111000001110000000111100000000011100000000000001111000000001110000001111100001111000000011110000000000000001110000111100000001111000001110000000011110000001111000000000000001110000001111100000000000000111110000001111000011110000000011110000001111000011111000000111100000111000011110000000000000011110000000111000000001110000000000000001110000011100000000000000000011110000000000001111000000111100000111000000111110000011100001111000000111110000111100000001111000000000000011100000;
  localparam words21  = 588'b000000011110000001111000011110000001111000011111100001111000000000000000001111000000000001111000111110000111111000001110000000111111100011111100000000000001111000000001111000011111100001111000000011110000000000000001110000111100000001111000001111111100001111000011110000000000000001111000011111100000000000000111111000011110000011110000000001111000011110000011111100001111000000111000001111100000111100011110000000111000000001110000000000000001110000011111111000000000000001111100001110000111100001111000000111100001111110000011100000111100001111110000111100000001111000000000000011111111;
  localparam words22  = 588'b000000011110000000111111111110000000111111111111100001111000000000000000001110000000000001111000111111111111110000001110000000011111111111111000000000000001111000000000111111111111100001111000000011110000000000000001110000111100000001111000001111111100000111111111110000000000000000111111111111100000000000000111111111111100000011110000000000111111111110000011111111111110000000111000000111111111111100011110000000111000000001110000000000000001110000011111111000000000000000111111111110000011111111111000000011111111111110000011100000011111111111110000111100000001111000000000000011111111;
  localparam words23  = 588'b000000011110000000011111111000000000011111110111100001111000000000000000011110000000000000111000011111111111100000001110000000000111111111110000000000000001111000000000011111110011100001111000000011110000000000000001110000111100000001111000000111111100000011111111000000000000000000011111110011100000000000000111101111111000000011110000000000011111111000000011110111111100000000111000000011111111111000011110000000111000000001110000000000000001110000001111111000000000000000011111111110000001111111100000000001111111011110000011100000001111111011110000111100000001111000000000000001111111;
  localparam words24  = 588'b000000000000000000000111100000000000000111000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000111110000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111000000000000000000000111100011100000000000000000000000000111100000000000000001110000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000011110000000000000011100000000000000000000000011100000000000000000000000000000000000000000000000;
  localparam words25  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words26  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words27  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words28  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words29  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words30  = 588'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words31  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words32  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words33  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words34  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words35  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words36  = 588'b001111000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words37  = 588'b001111001111100000000000111111100000000011000111110000000000001111100111100000111000000001111111000000000000000000001111111000000000110001111100000000000011111001111000000000000000110001111100000000000011111100000001110000000111000000011000000000000000110000111111111100000000000000110001111100000000000011111110000000000011111110000000000011111001111000000011111110000000000000001111111111000000011111100000000000000000001100011110000001111111000000000011111110000011111111110000001111111000000000110001111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words38  = 588'b001111011111111000000011111111111000000111101111111100000000111111111111100000111000000011111111100000000000000000111111111110000001111011111111000000001111111111111000000000000001111011111111000000001111111111000001110000001111000000111000000000000000111000111111111100000000000001111011111111000000000111111111000000000111111111000000001111111111111000001111111111100000000000001111111111000001111111111000000000000000011111111111000011111111100000001111111111100011111111110000111111111110000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words39  = 588'b001111111111111100000011111111111100000111111111111110000001111111111111100000111000000111111111110000000000000000111111111111000001111111111111100000011111111111111000000000000001111111111111100000011111111111100001111000001111100000111000000000000000111000111111111100000000000001111111111111100000001111111111100000001111111111100000011111111111111000011111111111100000000000001111111111000011111111111100000000000000011111111111000111111111110000011111111111100011111111110000111111111111000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words40  = 588'b001111110000111100000010000000111100000111111000011110000001111000011111100000111000001111000001111000000000000000100000001111000001111110000111100000011110000111111000000000000001111110000111100000011110000011110000111000001111100000111000000000000000111000011110000000000000000001111110000111100000011110000011110000011110000011110000011110000111111000011100000001000000000000000111100000000011110000011110000000000000011111100000001111000001111000011100000001000001111000000000100000001111000001111110000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words41  = 588'b001111100000011100000000000000011110000111110000001110000011110000001111100000111000011110000000111100000000000000000000000111100001111100000011100000111100000011111000000000000001111100000011100000111100000011110000111000011111100001111000000000000000111000011110000000000000000001111100000011100000111100000001111000111100000001111000111100000011111000011100000000000000000000000111100000000111100000011110000000000000011111000000011110000000111100011100000000000001111000000000000000000111100001111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words42  = 588'b001111000000011110000000000000001110000111100000001111000011100000000111100000111000011100000000011100000000000000000000000011100001111000000011110000111000000001111000000000000001111000000011110000111000000001111000111100011101100001110000000000000000111000011110000000000000000001111000000011110000111000000000111000111000000000111000111000000001111000111100000000000000000000000111100000000111000000001111000000000000011110000000011100000000011100111100000000000001111000000000000000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words43  = 588'b001111000000011110000000001111111110000111100000001111000011100000000111100000111000011100000000011100000000000000000011111111100001111000000011110000111000000001111000000000000001111000000011110000111000000001111000011100011101110001110000000000000000111000011110000000000000000001111000000011110000111000000000111000111000000000111000111000000001111000011110000000000000000000000111100000000111000000001111000000000000011110000000011100000000011100011110000000000001111000000000000011111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words44  = 588'b001111000000011110000001111111111110000111100000001111000111100000000111100000111000111111111111111100000000000000011111111111100001111000000011110001111000000001111000000000000001111000000011110001111000000001111000011100011101110011110000000000000000111000011110000000000000000001111000000011110001111111111111111001111111111111111001111000000001111000011111111000000000000000000111100000001111000000001111000000000000011110000000111111111111111100011111111000000001111000000000011111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words45  = 588'b001111000000011110000011111111111110000111100000001111000111100000000111100000111000111111111111111100000000000000111111111111100001111000000011110001111000000001111000000000000001111000000011110001111000000000111000011100111001110011100000000000000000111000011110000000000000000001111000000011110001111111111111111001111111111111111001111000000001111000001111111110000000000000000111100000001111000000000111000000000000011110000000111111111111111100001111111110000001111000000000111111111111100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words46  = 588'b001111000000011110000111100000001110000111100000001111000111100000000111100000111000111111111111111100000000000001111000000011100001111000000011110001111000000001111000000000000001111000000011110001111000000000111000011110111000110011100000000000000000111000011110000000000000000001111000000011110001111111111111111001111111111111111001111000000001111000000011111111000000000000000111100000001111000000000111000000000000011110000000111111111111111100000011111111000001111000000001111000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words47  = 588'b001111000000011110000111000000001110000111100000001111000111100000000111100000111000111100000000000000000000000001110000000011100001111000000011110001111000000001111000000000000001111000000011110001111000000001111000001110111000111011100000000000000000111000011110000000000000000001111000000011110001111000000000000001111000000000000001111000000001111000000000001111100000000000000111100000001111000000001111000000000000011110000000111100000000000000000000001111100001111000000001110000000011100001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words48  = 588'b001111000000011110000111000000011110000111100000001111000011100000000111100000111000011100000000000000000000000001110000000111100001111000000011110000111000000001111000000000000001111000000011110000111000000001111000001110110000111111100000000000000000111000001110000000000000000001111000000011110000111000000000000000111000000000000000111000000001111000000000000011100000000000000011100000000111000000001111000000000000011110000000011100000000000000000000000011100000111000000001110000000111100001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words49  = 588'b001111000000011110000111000000011110000111100000001111000011100000000111100000111000011110000000000000000000000001110000000111100001111000000011110000111000000001111000000000000001111000000011110000111100000001110000001111110000111111000000000000000000111000001110000000000000000001111000000011110000111100000000000000111100000000000000111000000001111000000000000011100000000000000011100000000111100000001110000000000000011110000000011110000000000000000000000011100000111000000001110000000111100001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000;
  localparam words50  = 588'b001111000000011110000111000000111110000111100000001111000011110000001111100000111000011110000000000000000000000001110000001111100001111000000011110000111100000011111000000000000001111000000011110000111100000011110000001111110000011111000000000000000000111000001110000000000000000001111000000011110000111100000000000000111100000000000000111100000011111000000000000011100000000000000011100000000111100000011110000000000000011110000000011110000000000000000000000011100000111000000001110000001111100001111000000000111000000000111000000000000000000000000000000000000000000000000000000000000000;
  localparam words51  = 588'b001111000000011110000111100001111110000111100000001111000001111000011111100000111000001111100000111100000000000001111000011111100001111000000011110000011110000111111000000000000001111000000011110000011110000111100000000111110000011111000000000000000000111000001111111100000000000001111000000011110000011111000001111000011111000001111000011110000111111000111100000111100000000000000011111111000011110000111100000000000000011110000000001111100000111100111100000111100000111111110001111000011111100001111000000000111111110000111100000000000000000000000000000000000000000000000000000000000000;
  localparam words52  = 588'b001111000000011110000011111111111110000111100000001111000000111111111111100000111000000111111111111100000000000000111111111111100001111000000011110000001111111111111000000000000001111000000011110000001111111111100000000111100000011111000000000000000000111000001111111100000000000001111000000011110000001111111111111000001111111111111000001111111111111000111111111111000000000000000011111111000001111111111100000000000000011110000000000111111111111100111111111111000000111111110000111111111111100001111000000000111111110000111100000000000000000000000000000000000000000000000000000000000000;
  localparam words53  = 588'b001111000000011110000001111111001110000111100000001111000000011111110111100000111000000011111111111000000000000000011111110011100001111000000011110000000111111101111000000000000001111000000011110000000111111110000000000111100000011110000000000000000000111000000111111100000000000001111000000011110000000111111111110000000111111111110000000111111101111000011111111110000000000000000001111111000000111111110000000000000000011110000000000011111111111000011111111110000000011111110000011111110011100001111000000000011111110000111100000000000000000000000000000000000000000000000000000000000000;
  localparam words54  = 588'b000000000000000000000000011100000000000000000000000000000000000111000000000000000000000000011111000000000000000000000111000000000000000000000000000000000001110000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000111110000000000001110000000000000011111000000000000000000000000000000000001111000000000000000000000000000000000000011111000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  wire            blank;
  reg             blank_h;
  reg             blank_v;

  assign blank = (blank_h | blank_v);

  // 2^10  = 1024
  reg [9:0]       count_h;
  // 2^15 = 32768
  reg [14:0]      count_v;

  wire            red;
  wire            grn;
  reg             blu;
  reg             wht;
  reg             hs_out;
  reg             vs_out;

  reg [3:0]       fb[3:0];

  assign r0 = red;
  assign r1 = red;
  assign r2 = red;
  assign r3 = red;
  assign b0 = blu;
  assign b1 = blu;
  assign b2 = blu;
  assign b3 = blu;
  assign g0 = grn;
  assign g1 = grn;
  assign g2 = grn;
  assign g3 = grn;
  assign hs = !hs_out;
  assign vs = !vs_out;

  assign red = wht;
  assign grn = wht;

  always @ (blank) begin
    if (blank) begin
      blu <= 1'b0;
      wht <= 1'b0;
    end else begin
      blu <= 1'b1;
      if (count_v > 99 && count_v < 212 && count_h > 79 && count_h < 139) begin
        case(count_v-99)
          1 : wht <= smile001[138-count_h];
          2 : wht <= smile002[138-count_h];
          3 : wht <= smile003[138-count_h];
          4 : wht <= smile004[138-count_h];
          5 : wht <= smile005[138-count_h];
          6 : wht <= smile006[138-count_h];
          7 : wht <= smile007[138-count_h];
          8 : wht <= smile008[138-count_h];
          9 : wht <= smile009[138-count_h];
          10 : wht <= smile010[138-count_h];
          11 : wht <= smile011[138-count_h];
          12 : wht <= smile012[138-count_h];
          13 : wht <= smile013[138-count_h];
          14 : wht <= smile014[138-count_h];
          15 : wht <= smile015[138-count_h];
          16 : wht <= smile016[138-count_h];
          17 : wht <= smile017[138-count_h];
          18 : wht <= smile018[138-count_h];
          19 : wht <= smile019[138-count_h];
          20 : wht <= smile020[138-count_h];
          21 : wht <= smile021[138-count_h];
          22 : wht <= smile022[138-count_h];
          23 : wht <= smile023[138-count_h];
          24 : wht <= smile024[138-count_h];
          25 : wht <= smile025[138-count_h];
          26 : wht <= smile026[138-count_h];
          27 : wht <= smile027[138-count_h];
          28 : wht <= smile028[138-count_h];
          29 : wht <= smile029[138-count_h];
          30 : wht <= smile030[138-count_h];
          31 : wht <= smile031[138-count_h];
          32 : wht <= smile032[138-count_h];
          33 : wht <= smile033[138-count_h];
          34 : wht <= smile034[138-count_h];
          35 : wht <= smile035[138-count_h];
          36 : wht <= smile036[138-count_h];
          37 : wht <= smile037[138-count_h];
          38 : wht <= smile038[138-count_h];
          39 : wht <= smile039[138-count_h];
          40 : wht <= smile040[138-count_h];
          41 : wht <= smile041[138-count_h];
          42 : wht <= smile042[138-count_h];
          43 : wht <= smile043[138-count_h];
          44 : wht <= smile044[138-count_h];
          45 : wht <= smile045[138-count_h];
          46 : wht <= smile046[138-count_h];
          47 : wht <= smile047[138-count_h];
          48 : wht <= smile048[138-count_h];
          49 : wht <= smile049[138-count_h];
          50 : wht <= smile050[138-count_h];
          51 : wht <= smile051[138-count_h];
          52 : wht <= smile052[138-count_h];
          53 : wht <= smile053[138-count_h];
          54 : wht <= smile054[138-count_h];
          55 : wht <= smile055[138-count_h];
          56 : wht <= smile056[138-count_h];
          57 : wht <= smile057[138-count_h];
          58 : wht <= smile058[138-count_h];
          59 : wht <= smile059[138-count_h];
          60 : wht <= smile060[138-count_h];
          61 : wht <= smile061[138-count_h];
          62 : wht <= smile062[138-count_h];
          63 : wht <= smile063[138-count_h];
          64 : wht <= smile064[138-count_h];
          65 : wht <= smile065[138-count_h];
          66 : wht <= smile066[138-count_h];
          67 : wht <= smile067[138-count_h];
          68 : wht <= smile068[138-count_h];
          69 : wht <= smile069[138-count_h];
          70 : wht <= smile070[138-count_h];
          71 : wht <= smile071[138-count_h];
          72 : wht <= smile072[138-count_h];
          73 : wht <= smile073[138-count_h];
          74 : wht <= smile074[138-count_h];
          75 : wht <= smile075[138-count_h];
          76 : wht <= smile076[138-count_h];
          77 : wht <= smile077[138-count_h];
          78 : wht <= smile078[138-count_h];
          79 : wht <= smile079[138-count_h];
          80 : wht <= smile080[138-count_h];
          81 : wht <= smile081[138-count_h];
          82 : wht <= smile082[138-count_h];
          83 : wht <= smile083[138-count_h];
          84 : wht <= smile084[138-count_h];
          85 : wht <= smile085[138-count_h];
          86 : wht <= smile086[138-count_h];
          87 : wht <= smile087[138-count_h];
          88 : wht <= smile088[138-count_h];
          89 : wht <= smile089[138-count_h];
          90 : wht <= smile090[138-count_h];
          91 : wht <= smile091[138-count_h];
          92 : wht <= smile092[138-count_h];
          93 : wht <= smile093[138-count_h];
          94 : wht <= smile094[138-count_h];
          95 : wht <= smile095[138-count_h];
          96 : wht <= smile096[138-count_h];
          97 : wht <= smile097[138-count_h];
          98 : wht <= smile098[138-count_h];
          99 : wht <= smile099[138-count_h];
          100 : wht <= smile100[138-count_h];
          101 : wht <= smile101[138-count_h];
          102 : wht <= smile102[138-count_h];
          103 : wht <= smile103[138-count_h];
          104 : wht <= smile104[138-count_h];
          105 : wht <= smile105[138-count_h];
          106 : wht <= smile106[138-count_h];
          107 : wht <= smile107[138-count_h];
          108 : wht <= smile108[138-count_h];
          109 : wht <= smile109[138-count_h];
          110 : wht <= smile110[138-count_h];
          111 : wht <= smile111[138-count_h];
          112 : wht <= smile112[138-count_h];
          default: wht <= 1'b0;
        endcase
//       end else if (count_v > 299 && count_v < 354 && count_h > 14 && count_h < 602) begin
//         case(count_v-299)
//           1 : wht  <= words01[602-count_h];
//           2 : wht  <= words02[602-count_h];
//           3 : wht  <= words03[602-count_h];
//           4 : wht  <= words04[602-count_h];
//           5 : wht  <= words05[602-count_h];
//           6 : wht  <= words06[602-count_h];
//           7 : wht  <= words07[602-count_h];
//           8 : wht  <= words08[602-count_h];
//           9 : wht  <= words09[602-count_h];
//           10 : wht <= words10[602-count_h];
//           11 : wht <= words11[602-count_h];
//           12 : wht <= words12[602-count_h];
//           13 : wht <= words13[602-count_h];
//           14 : wht <= words14[602-count_h];
//           15 : wht <= words15[602-count_h];
//           16 : wht <= words16[602-count_h];
//           17 : wht <= words17[602-count_h];
//           18 : wht <= words18[602-count_h];
//           19 : wht <= words19[602-count_h];
//           20 : wht <= words20[602-count_h];
//           21 : wht <= words21[602-count_h];
//           22 : wht <= words22[602-count_h];
//           23 : wht <= words23[602-count_h];
//           24 : wht <= words24[602-count_h];
//           25 : wht <= words25[602-count_h];
//           26 : wht <= words26[602-count_h];
//           27 : wht <= words27[602-count_h];
//           28 : wht <= words28[602-count_h];
//           29 : wht <= words29[602-count_h];
//           30 : wht <= words30[602-count_h];
//           31 : wht <= words31[602-count_h];
//           32 : wht <= words32[602-count_h];
//           33 : wht <= words33[602-count_h];
//           34 : wht <= words34[602-count_h];
//           35 : wht <= words35[602-count_h];
//           36 : wht <= words36[602-count_h];
//           37 : wht <= words37[602-count_h];
//           38 : wht <= words38[602-count_h];
//           39 : wht <= words39[602-count_h];
//           40 : wht <= words40[602-count_h];
//           41 : wht <= words41[602-count_h];
//           42 : wht <= words42[602-count_h];
//           43 : wht <= words43[602-count_h];
//           44 : wht <= words44[602-count_h];
//           45 : wht <= words45[602-count_h];
//           46 : wht <= words46[602-count_h];
//           47 : wht <= words47[602-count_h];
//           48 : wht <= words48[602-count_h];
//           49 : wht <= words49[602-count_h];
//           50 : wht <= words50[602-count_h];
//           51 : wht <= words51[602-count_h];
//           52 : wht <= words52[602-count_h];
//           53 : wht <= words53[602-count_h];
//           54 : wht <= words54[602-count_h];
//           default: wht <= 1'b0;
//         endcase
      end else begin
        wht <= 1'b0;
      end
    end
  end

  always @ (posedge clk) begin
    hs_out <= 1'b0;
    if (rst) begin
      count_h <= 10'b11_1111_1111;
      blank_h <= 1'b1;
    end else if (count_h < h_visible) begin
	  // horizontal visible
      count_h <= count_h + 1;
    end else if (count_h < h_frontporch) begin
	  // horizontal front porch
      count_h <= count_h + 1;
      blank_h <= 1'b1;
    end else if (count_h < h_sync) begin
	  // horizontal sync
      count_h <= count_h + 1;
	  hs_out <= 1'b1;
    end else if (count_h < h_backporch) begin
	  // horizontal back porch
      count_h <= count_h + 1;
    end else begin
      count_h <= 1;
      blank_h <= 1'b0;
    end
  end

  always @ (posedge clk) begin
    if (rst) begin
      count_v <= 15'b111_1111_1111_1111;
      blank_v <= 1'b1;
      vs_out  <= 1'b0;
    end else if (count_h >= h_backporch) begin
      if (count_v < v_visible) begin
        count_v <= count_v + 1;
      end else if (count_v < v_backporch) begin
        count_v <= count_v + 1;
        blank_v <= 1'b1;
        if (count_v > v_frontporch && count_v < v_sync) begin
          vs_out <= 1'b1;
        end else begin
          vs_out <= 1'b0;
        end
      end else begin
        count_v <= 1;
        blank_v <= 1'b0;
      end
    end
  end
  
endmodule
